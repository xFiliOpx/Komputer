<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-136.173,297.585,133.88,93.2654</PageViewport>
<gate>
<ID>389</ID>
<type>AA_AND2</type>
<position>-66.5,277</position>
<input>
<ID>IN_0</ID>375 </input>
<input>
<ID>IN_1</ID>366 </input>
<output>
<ID>OUT</ID>358 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1</ID>
<type>AE_DFF_LOW</type>
<position>12.5,210.5</position>
<input>
<ID>IN_0</ID>14 </input>
<output>
<ID>OUT_0</ID>9 </output>
<input>
<ID>clock</ID>13 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>2</ID>
<type>AE_DFF_LOW</type>
<position>21.5,210.5</position>
<input>
<ID>IN_0</ID>9 </input>
<output>
<ID>OUT_0</ID>10 </output>
<input>
<ID>clock</ID>13 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3</ID>
<type>AE_DFF_LOW</type>
<position>30.5,210.5</position>
<input>
<ID>IN_0</ID>10 </input>
<output>
<ID>OUT_0</ID>12 </output>
<input>
<ID>clock</ID>13 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>393</ID>
<type>AE_SMALL_INVERTER</type>
<position>37,230.5</position>
<input>
<ID>IN_0</ID>11 </input>
<output>
<ID>OUT_0</ID>375 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5</ID>
<type>AE_OR2</type>
<position>37,225</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>9</ID>
<type>BE_ROM_8x8</type>
<position>-37.5,251.5</position>
<input>
<ID>ADDRESS_0</ID>38 </input>
<input>
<ID>ADDRESS_1</ID>29 </input>
<input>
<ID>ADDRESS_2</ID>32 </input>
<input>
<ID>ADDRESS_3</ID>37 </input>
<input>
<ID>ADDRESS_4</ID>30 </input>
<input>
<ID>ADDRESS_5</ID>35 </input>
<input>
<ID>ADDRESS_6</ID>31 </input>
<input>
<ID>ADDRESS_7</ID>33 </input>
<output>
<ID>DATA_OUT_0</ID>24 </output>
<output>
<ID>DATA_OUT_1</ID>25 </output>
<output>
<ID>DATA_OUT_2</ID>23 </output>
<output>
<ID>DATA_OUT_3</ID>28 </output>
<output>
<ID>DATA_OUT_4</ID>27 </output>
<output>
<ID>DATA_OUT_5</ID>26 </output>
<output>
<ID>DATA_OUT_6</ID>34 </output>
<output>
<ID>DATA_OUT_7</ID>36 </output>
<input>
<ID>ENABLE_0</ID>40 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam>
<lparam>Address:7 2</lparam>
<lparam>Address:8 5</lparam>
<lparam>Address:29 2</lparam>
<lparam>Address:30 255</lparam></gate>
<gate>
<ID>11</ID>
<type>HA_JUNC_2</type>
<position>-43.5,248</position>
<input>
<ID>N_in0</ID>15 </input>
<input>
<ID>N_in1</ID>38 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>HA_JUNC_2</type>
<position>-43.5,249</position>
<input>
<ID>N_in0</ID>16 </input>
<input>
<ID>N_in1</ID>29 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>13</ID>
<type>HA_JUNC_2</type>
<position>-43.5,250</position>
<input>
<ID>N_in0</ID>17 </input>
<input>
<ID>N_in1</ID>32 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>HA_JUNC_2</type>
<position>-43.5,251</position>
<input>
<ID>N_in0</ID>18 </input>
<input>
<ID>N_in1</ID>37 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>HA_JUNC_2</type>
<position>-43.5,252</position>
<input>
<ID>N_in0</ID>19 </input>
<input>
<ID>N_in1</ID>30 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>HA_JUNC_2</type>
<position>-43.5,253</position>
<input>
<ID>N_in0</ID>20 </input>
<input>
<ID>N_in1</ID>35 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>17</ID>
<type>HA_JUNC_2</type>
<position>-43.5,254</position>
<input>
<ID>N_in0</ID>21 </input>
<input>
<ID>N_in1</ID>31 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>HA_JUNC_2</type>
<position>-43.5,255</position>
<input>
<ID>N_in0</ID>22 </input>
<input>
<ID>N_in1</ID>33 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>408</ID>
<type>BE_NOR2</type>
<position>30,309.5</position>
<input>
<ID>IN_0</ID>391 </input>
<input>
<ID>IN_1</ID>388 </input>
<output>
<ID>OUT</ID>387 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>20</ID>
<type>HA_JUNC_2</type>
<position>-41,243.5</position>
<input>
<ID>N_in0</ID>62 </input>
<input>
<ID>N_in1</ID>36 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>409</ID>
<type>BE_NOR2</type>
<position>34,309.5</position>
<input>
<ID>IN_0</ID>387 </input>
<input>
<ID>IN_1</ID>392 </input>
<output>
<ID>OUT</ID>388 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>21</ID>
<type>HA_JUNC_2</type>
<position>-40,243.5</position>
<input>
<ID>N_in0</ID>61 </input>
<input>
<ID>N_in1</ID>34 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>22</ID>
<type>HA_JUNC_2</type>
<position>-39,243.5</position>
<input>
<ID>N_in0</ID>60 </input>
<input>
<ID>N_in1</ID>26 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>23</ID>
<type>HA_JUNC_2</type>
<position>-38,243.5</position>
<input>
<ID>N_in0</ID>59 </input>
<input>
<ID>N_in1</ID>27 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>24</ID>
<type>HA_JUNC_2</type>
<position>-37,243.5</position>
<input>
<ID>N_in0</ID>58 </input>
<input>
<ID>N_in1</ID>28 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>25</ID>
<type>HA_JUNC_2</type>
<position>-36,243.5</position>
<input>
<ID>N_in0</ID>57 </input>
<input>
<ID>N_in1</ID>23 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>26</ID>
<type>HA_JUNC_2</type>
<position>-35,243.5</position>
<input>
<ID>N_in0</ID>56 </input>
<input>
<ID>N_in1</ID>25 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>27</ID>
<type>HA_JUNC_2</type>
<position>-34,243.5</position>
<input>
<ID>N_in0</ID>55 </input>
<input>
<ID>N_in1</ID>24 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>417</ID>
<type>HA_JUNC_2</type>
<position>30,314</position>
<input>
<ID>N_in0</ID>387 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>419</ID>
<type>HA_JUNC_2</type>
<position>34,314</position>
<input>
<ID>N_in0</ID>388 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>31</ID>
<type>EE_VDD</type>
<position>-31.5,252</position>
<output>
<ID>OUT_0</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>420</ID>
<type>HA_JUNC_2</type>
<position>30,305</position>
<input>
<ID>N_in0</ID>393 </input>
<input>
<ID>N_in1</ID>391 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>32</ID>
<type>HA_JUNC_2</type>
<position>-32,210.5</position>
<input>
<ID>N_in0</ID>57 </input>
<input>
<ID>N_in1</ID>42 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>421</ID>
<type>HA_JUNC_2</type>
<position>34,305</position>
<input>
<ID>N_in0</ID>394 </input>
<input>
<ID>N_in1</ID>392 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>33</ID>
<type>HA_JUNC_2</type>
<position>-32,214.5</position>
<input>
<ID>N_in0</ID>55 </input>
<input>
<ID>N_in1</ID>41 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>423</ID>
<type>AA_TOGGLE</type>
<position>30,301.5</position>
<output>
<ID>OUT_0</ID>393 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>425</ID>
<type>AA_TOGGLE</type>
<position>34,301.5</position>
<output>
<ID>OUT_0</ID>394 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>37</ID>
<type>HA_JUNC_2</type>
<position>-32,208.5</position>
<input>
<ID>N_in0</ID>58 </input>
<input>
<ID>N_in1</ID>43 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>426</ID>
<type>BE_NOR2</type>
<position>-31,238.5</position>
<input>
<ID>IN_0</ID>397 </input>
<input>
<ID>IN_1</ID>396 </input>
<output>
<ID>OUT</ID>395 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>38</ID>
<type>HA_JUNC_2</type>
<position>-32,206.5</position>
<input>
<ID>N_in0</ID>59 </input>
<input>
<ID>N_in1</ID>44 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>427</ID>
<type>BE_NOR2</type>
<position>-27,238.5</position>
<input>
<ID>IN_0</ID>395 </input>
<input>
<ID>IN_1</ID>398 </input>
<output>
<ID>OUT</ID>396 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>39</ID>
<type>HA_JUNC_2</type>
<position>-32,204.5</position>
<input>
<ID>N_in0</ID>60 </input>
<input>
<ID>N_in1</ID>45 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>428</ID>
<type>HA_JUNC_2</type>
<position>-31,243</position>
<input>
<ID>N_in0</ID>395 </input>
<input>
<ID>N_in1</ID>1 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>40</ID>
<type>HA_JUNC_2</type>
<position>-32,202.5</position>
<input>
<ID>N_in0</ID>61 </input>
<input>
<ID>N_in1</ID>46 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>HA_JUNC_2</type>
<position>-32,200.5</position>
<input>
<ID>N_in0</ID>62 </input>
<input>
<ID>N_in1</ID>48 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>430</ID>
<type>HA_JUNC_2</type>
<position>-31,234</position>
<input>
<ID>N_in0</ID>12 </input>
<input>
<ID>N_in1</ID>397 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>431</ID>
<type>HA_JUNC_2</type>
<position>-27,234</position>
<input>
<ID>N_in0</ID>456 </input>
<input>
<ID>N_in1</ID>398 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>432</ID>
<type>BE_NOR2</type>
<position>-22.5,239</position>
<input>
<ID>IN_0</ID>409 </input>
<input>
<ID>IN_1</ID>408 </input>
<output>
<ID>OUT</ID>407 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>433</ID>
<type>BE_NOR2</type>
<position>-18.5,239</position>
<input>
<ID>IN_0</ID>407 </input>
<input>
<ID>IN_1</ID>410 </input>
<output>
<ID>OUT</ID>408 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>434</ID>
<type>HA_JUNC_2</type>
<position>-22.5,243.5</position>
<input>
<ID>N_in0</ID>407 </input>
<input>
<ID>N_in1</ID>2 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>435</ID>
<type>HA_JUNC_2</type>
<position>-22.5,234.5</position>
<input>
<ID>N_in0</ID>12 </input>
<input>
<ID>N_in1</ID>409 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>436</ID>
<type>HA_JUNC_2</type>
<position>-18.5,234.5</position>
<input>
<ID>N_in0</ID>457 </input>
<input>
<ID>N_in1</ID>410 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>48</ID>
<type>DA_FROM</type>
<position>11.5,205.5</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>437</ID>
<type>BE_NOR2</type>
<position>-14,239.5</position>
<input>
<ID>IN_0</ID>415 </input>
<input>
<ID>IN_1</ID>414 </input>
<output>
<ID>OUT</ID>413 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>438</ID>
<type>BE_NOR2</type>
<position>-10,239.5</position>
<input>
<ID>IN_0</ID>413 </input>
<input>
<ID>IN_1</ID>416 </input>
<output>
<ID>OUT</ID>414 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_AND2</type>
<position>-16,213.5</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>81 </input>
<output>
<ID>OUT</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>439</ID>
<type>HA_JUNC_2</type>
<position>-14,244</position>
<input>
<ID>N_in0</ID>413 </input>
<input>
<ID>N_in1</ID>3 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>51</ID>
<type>AA_AND2</type>
<position>-16,209.5</position>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>81 </input>
<output>
<ID>OUT</ID>73 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>440</ID>
<type>HA_JUNC_2</type>
<position>-14,235</position>
<input>
<ID>N_in0</ID>12 </input>
<input>
<ID>N_in1</ID>415 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>52</ID>
<type>AA_AND2</type>
<position>-16,205.5</position>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>81 </input>
<output>
<ID>OUT</ID>66 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>441</ID>
<type>HA_JUNC_2</type>
<position>-10,235</position>
<input>
<ID>N_in0</ID>458 </input>
<input>
<ID>N_in1</ID>416 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>53</ID>
<type>AA_AND2</type>
<position>-16,201.5</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>IN_1</ID>81 </input>
<output>
<ID>OUT</ID>65 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>442</ID>
<type>BE_NOR2</type>
<position>-5.5,240</position>
<input>
<ID>IN_0</ID>420 </input>
<input>
<ID>IN_1</ID>419 </input>
<output>
<ID>OUT</ID>418 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>443</ID>
<type>BE_NOR2</type>
<position>-1.5,240</position>
<input>
<ID>IN_0</ID>418 </input>
<input>
<ID>IN_1</ID>421 </input>
<output>
<ID>OUT</ID>419 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>55</ID>
<type>AE_OR3</type>
<position>-1,199</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>10 </input>
<input>
<ID>IN_2</ID>9 </input>
<output>
<ID>OUT</ID>80 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>444</ID>
<type>HA_JUNC_2</type>
<position>-5.5,244.5</position>
<input>
<ID>N_in0</ID>418 </input>
<input>
<ID>N_in1</ID>4 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>445</ID>
<type>HA_JUNC_2</type>
<position>-5.5,235.5</position>
<input>
<ID>N_in0</ID>12 </input>
<input>
<ID>N_in1</ID>420 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>57</ID>
<type>AE_SMALL_INVERTER</type>
<position>-10,213.5</position>
<input>
<ID>IN_0</ID>64 </input>
<output>
<ID>OUT_0</ID>72 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>446</ID>
<type>HA_JUNC_2</type>
<position>-1.5,235.5</position>
<input>
<ID>N_in0</ID>459 </input>
<input>
<ID>N_in1</ID>421 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>58</ID>
<type>AE_SMALL_INVERTER</type>
<position>-10,205.5</position>
<input>
<ID>IN_0</ID>66 </input>
<output>
<ID>OUT_0</ID>74 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>447</ID>
<type>BE_NOR2</type>
<position>3,240.5</position>
<input>
<ID>IN_0</ID>425 </input>
<input>
<ID>IN_1</ID>424 </input>
<output>
<ID>OUT</ID>423 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>59</ID>
<type>AE_SMALL_INVERTER</type>
<position>-10,201.5</position>
<input>
<ID>IN_0</ID>65 </input>
<output>
<ID>OUT_0</ID>75 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>448</ID>
<type>BE_NOR2</type>
<position>7,240.5</position>
<input>
<ID>IN_0</ID>423 </input>
<input>
<ID>IN_1</ID>426 </input>
<output>
<ID>OUT</ID>424 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>60</ID>
<type>AA_AND2</type>
<position>-16,196.5</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>81 </input>
<output>
<ID>OUT</ID>67 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>449</ID>
<type>HA_JUNC_2</type>
<position>3,245</position>
<input>
<ID>N_in0</ID>423 </input>
<input>
<ID>N_in1</ID>5 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>61</ID>
<type>AA_AND2</type>
<position>-16,192.5</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>81 </input>
<output>
<ID>OUT</ID>70 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>450</ID>
<type>HA_JUNC_2</type>
<position>3,236</position>
<input>
<ID>N_in0</ID>12 </input>
<input>
<ID>N_in1</ID>425 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>62</ID>
<type>AA_AND2</type>
<position>-16,188.5</position>
<input>
<ID>IN_0</ID>46 </input>
<input>
<ID>IN_1</ID>81 </input>
<output>
<ID>OUT</ID>69 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>451</ID>
<type>HA_JUNC_2</type>
<position>7,236</position>
<input>
<ID>N_in0</ID>460 </input>
<input>
<ID>N_in1</ID>426 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>63</ID>
<type>AA_AND2</type>
<position>-16,184.5</position>
<input>
<ID>IN_0</ID>48 </input>
<input>
<ID>IN_1</ID>81 </input>
<output>
<ID>OUT</ID>68 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>452</ID>
<type>BE_NOR2</type>
<position>11.5,241</position>
<input>
<ID>IN_0</ID>429 </input>
<input>
<ID>IN_1</ID>428 </input>
<output>
<ID>OUT</ID>427 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>64</ID>
<type>AE_SMALL_INVERTER</type>
<position>-10,196.5</position>
<input>
<ID>IN_0</ID>67 </input>
<output>
<ID>OUT_0</ID>76 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>453</ID>
<type>BE_NOR2</type>
<position>15.5,241</position>
<input>
<ID>IN_0</ID>427 </input>
<input>
<ID>IN_1</ID>430 </input>
<output>
<ID>OUT</ID>428 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>65</ID>
<type>AE_SMALL_INVERTER</type>
<position>-10,188.5</position>
<input>
<ID>IN_0</ID>69 </input>
<output>
<ID>OUT_0</ID>78 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>454</ID>
<type>HA_JUNC_2</type>
<position>11.5,245.5</position>
<input>
<ID>N_in0</ID>427 </input>
<input>
<ID>N_in1</ID>6 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>66</ID>
<type>AE_SMALL_INVERTER</type>
<position>-10,184.5</position>
<input>
<ID>IN_0</ID>68 </input>
<output>
<ID>OUT_0</ID>77 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>455</ID>
<type>HA_JUNC_2</type>
<position>11.5,236.5</position>
<input>
<ID>N_in0</ID>12 </input>
<input>
<ID>N_in1</ID>429 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>67</ID>
<type>AE_SMALL_INVERTER</type>
<position>-10,192.5</position>
<input>
<ID>IN_0</ID>70 </input>
<output>
<ID>OUT_0</ID>79 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>456</ID>
<type>HA_JUNC_2</type>
<position>15.5,236.5</position>
<input>
<ID>N_in0</ID>461 </input>
<input>
<ID>N_in1</ID>430 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>457</ID>
<type>BE_NOR2</type>
<position>20,241.5</position>
<input>
<ID>IN_0</ID>433 </input>
<input>
<ID>IN_1</ID>432 </input>
<output>
<ID>OUT</ID>431 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>69</ID>
<type>AE_SMALL_INVERTER</type>
<position>-9,199</position>
<input>
<ID>IN_0</ID>80 </input>
<output>
<ID>OUT_0</ID>81 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>458</ID>
<type>BE_NOR2</type>
<position>24,241.5</position>
<input>
<ID>IN_0</ID>431 </input>
<input>
<ID>IN_1</ID>434 </input>
<output>
<ID>OUT</ID>432 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>459</ID>
<type>HA_JUNC_2</type>
<position>20,246</position>
<input>
<ID>N_in0</ID>431 </input>
<input>
<ID>N_in1</ID>7 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>460</ID>
<type>HA_JUNC_2</type>
<position>20,237</position>
<input>
<ID>N_in0</ID>12 </input>
<input>
<ID>N_in1</ID>433 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>461</ID>
<type>HA_JUNC_2</type>
<position>24,237</position>
<input>
<ID>N_in0</ID>462 </input>
<input>
<ID>N_in1</ID>434 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>462</ID>
<type>BE_NOR2</type>
<position>28.5,242</position>
<input>
<ID>IN_0</ID>437 </input>
<input>
<ID>IN_1</ID>436 </input>
<output>
<ID>OUT</ID>435 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>463</ID>
<type>BE_NOR2</type>
<position>32.5,242</position>
<input>
<ID>IN_0</ID>435 </input>
<input>
<ID>IN_1</ID>438 </input>
<output>
<ID>OUT</ID>436 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>464</ID>
<type>HA_JUNC_2</type>
<position>28.5,246.5</position>
<input>
<ID>N_in0</ID>435 </input>
<input>
<ID>N_in1</ID>8 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>465</ID>
<type>HA_JUNC_2</type>
<position>28.5,237.5</position>
<input>
<ID>N_in0</ID>12 </input>
<input>
<ID>N_in1</ID>437 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>466</ID>
<type>HA_JUNC_2</type>
<position>32.5,237.5</position>
<input>
<ID>N_in0</ID>463 </input>
<input>
<ID>N_in1</ID>438 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>468</ID>
<type>AA_AND2</type>
<position>-27,229.5</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>456 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>469</ID>
<type>AA_AND2</type>
<position>-18.5,230</position>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>457 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>470</ID>
<type>AA_AND2</type>
<position>-10,230.5</position>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>458 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>471</ID>
<type>AA_AND2</type>
<position>-1.5,231</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>459 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>472</ID>
<type>AA_AND2</type>
<position>7,231.5</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>460 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>473</ID>
<type>AA_AND2</type>
<position>15.5,232</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>461 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>474</ID>
<type>AA_AND2</type>
<position>24,232.5</position>
<input>
<ID>IN_0</ID>46 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>462 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>475</ID>
<type>AA_AND2</type>
<position>32.5,233</position>
<input>
<ID>IN_0</ID>48 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>463 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>179</ID>
<type>AA_RAM_4x4</type>
<position>38.5,150.5</position>
<input>
<ID>ADDRESS_0</ID>205 </input>
<input>
<ID>ADDRESS_1</ID>203 </input>
<input>
<ID>ADDRESS_2</ID>202 </input>
<input>
<ID>ADDRESS_3</ID>204 </input>
<input>
<ID>DATA_IN_0</ID>213 </input>
<input>
<ID>DATA_IN_1</ID>214 </input>
<input>
<ID>DATA_IN_2</ID>216 </input>
<input>
<ID>DATA_IN_3</ID>215 </input>
<output>
<ID>DATA_OUT_0</ID>213 </output>
<output>
<ID>DATA_OUT_1</ID>214 </output>
<output>
<ID>DATA_OUT_2</ID>216 </output>
<output>
<ID>DATA_OUT_3</ID>215 </output>
<input>
<ID>ENABLE_0</ID>218 </input>
<input>
<ID>write_clock</ID>219 </input>
<input>
<ID>write_enable</ID>227 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 4</lparam>
<lparam>DATA_BITS 4</lparam>
<lparam>Address:0 2</lparam>
<lparam>Address:2 2</lparam>
<lparam>Address:6 11</lparam></gate>
<gate>
<ID>183</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>60,133.5</position>
<input>
<ID>IN_0</ID>224 </input>
<input>
<ID>IN_1</ID>223 </input>
<input>
<ID>IN_2</ID>225 </input>
<input>
<ID>IN_3</ID>226 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>185</ID>
<type>DD_KEYPAD_HEX</type>
<position>24,152</position>
<output>
<ID>OUT_0</ID>205 </output>
<output>
<ID>OUT_1</ID>203 </output>
<output>
<ID>OUT_2</ID>202 </output>
<output>
<ID>OUT_3</ID>204 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>201</ID>
<type>DD_KEYPAD_HEX</type>
<position>10.5,129.5</position>
<output>
<ID>OUT_0</ID>250 </output>
<output>
<ID>OUT_1</ID>233 </output>
<output>
<ID>OUT_2</ID>232 </output>
<output>
<ID>OUT_3</ID>228 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 2</lparam></gate>
<gate>
<ID>203</ID>
<type>AA_AND2</type>
<position>35,139.5</position>
<input>
<ID>IN_0</ID>227 </input>
<input>
<ID>IN_1</ID>250 </input>
<output>
<ID>OUT</ID>213 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>205</ID>
<type>AA_AND2</type>
<position>31,139.5</position>
<input>
<ID>IN_0</ID>227 </input>
<input>
<ID>IN_1</ID>233 </input>
<output>
<ID>OUT</ID>214 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>206</ID>
<type>AA_AND2</type>
<position>27,139.5</position>
<input>
<ID>IN_0</ID>227 </input>
<input>
<ID>IN_1</ID>232 </input>
<output>
<ID>OUT</ID>216 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>207</ID>
<type>AA_AND2</type>
<position>23,139.5</position>
<input>
<ID>IN_0</ID>227 </input>
<input>
<ID>IN_1</ID>228 </input>
<output>
<ID>OUT</ID>215 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>211</ID>
<type>AA_AND2</type>
<position>43,139.5</position>
<input>
<ID>IN_0</ID>218 </input>
<input>
<ID>IN_1</ID>215 </input>
<output>
<ID>OUT</ID>226 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>212</ID>
<type>AA_AND2</type>
<position>47,139.5</position>
<input>
<ID>IN_0</ID>218 </input>
<input>
<ID>IN_1</ID>216 </input>
<output>
<ID>OUT</ID>225 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>213</ID>
<type>AA_AND2</type>
<position>51,139.5</position>
<input>
<ID>IN_0</ID>218 </input>
<input>
<ID>IN_1</ID>214 </input>
<output>
<ID>OUT</ID>223 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>214</ID>
<type>AA_AND2</type>
<position>55,139.5</position>
<input>
<ID>IN_0</ID>218 </input>
<input>
<ID>IN_1</ID>213 </input>
<output>
<ID>OUT</ID>224 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>216</ID>
<type>AA_TOGGLE</type>
<position>58,150</position>
<output>
<ID>OUT_0</ID>218 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>218</ID>
<type>BB_CLOCK</type>
<position>38.5,156.5</position>
<output>
<ID>CLK</ID>219 </output>
<gparam>angle 0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>220</ID>
<type>AA_TOGGLE</type>
<position>54.5,151</position>
<output>
<ID>OUT_0</ID>227 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>268</ID>
<type>BB_CLOCK</type>
<position>-1,268.5</position>
<output>
<ID>CLK</ID>302 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 10</lparam></gate>
<gate>
<ID>270</ID>
<type>AE_SMALL_INVERTER</type>
<position>6.5,269.5</position>
<input>
<ID>IN_0</ID>302 </input>
<output>
<ID>OUT_0</ID>301 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>272</ID>
<type>DE_TO</type>
<position>11,269.5</position>
<input>
<ID>IN_0</ID>301 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID nclk</lparam></gate>
<gate>
<ID>274</ID>
<type>DE_TO</type>
<position>11,267.5</position>
<input>
<ID>IN_0</ID>302 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>290</ID>
<type>AE_DFF_LOW</type>
<position>-67,237</position>
<input>
<ID>IN_0</ID>231 </input>
<output>
<ID>OUT_0</ID>242 </output>
<input>
<ID>clock</ID>264 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>291</ID>
<type>AE_DFF_LOW</type>
<position>-67,228</position>
<input>
<ID>IN_0</ID>234 </input>
<output>
<ID>OUT_0</ID>243 </output>
<input>
<ID>clock</ID>264 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>293</ID>
<type>AE_DFF_LOW</type>
<position>-67,246</position>
<input>
<ID>IN_0</ID>230 </input>
<output>
<ID>OUT_0</ID>241 </output>
<input>
<ID>clock</ID>264 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>294</ID>
<type>AE_DFF_LOW</type>
<position>-67,219</position>
<input>
<ID>IN_0</ID>235 </input>
<output>
<ID>OUT_0</ID>244 </output>
<input>
<ID>clock</ID>264 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>296</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-72.5,255</position>
<input>
<ID>IN_0</ID>334 </input>
<input>
<ID>IN_1</ID>335 </input>
<input>
<ID>IN_2</ID>336 </input>
<input>
<ID>IN_3</ID>337 </input>
<input>
<ID>IN_B_0</ID>240 </input>
<output>
<ID>OUT_0</ID>230 </output>
<output>
<ID>OUT_1</ID>231 </output>
<output>
<ID>OUT_2</ID>234 </output>
<output>
<ID>OUT_3</ID>235 </output>
<output>
<ID>carry_out</ID>229 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>298</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-89.5,255</position>
<input>
<ID>IN_0</ID>333 </input>
<input>
<ID>IN_1</ID>338 </input>
<input>
<ID>IN_2</ID>339 </input>
<input>
<ID>IN_3</ID>340 </input>
<output>
<ID>OUT_0</ID>236 </output>
<output>
<ID>OUT_1</ID>237 </output>
<output>
<ID>OUT_2</ID>238 </output>
<output>
<ID>OUT_3</ID>239 </output>
<input>
<ID>carry_in</ID>229 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>299</ID>
<type>AE_DFF_LOW</type>
<position>-67,201</position>
<input>
<ID>IN_0</ID>237 </input>
<output>
<ID>OUT_0</ID>246 </output>
<input>
<ID>clock</ID>264 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>300</ID>
<type>AE_DFF_LOW</type>
<position>-67,192</position>
<input>
<ID>IN_0</ID>238 </input>
<output>
<ID>OUT_0</ID>247 </output>
<input>
<ID>clock</ID>264 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>301</ID>
<type>AE_DFF_LOW</type>
<position>-67,210</position>
<input>
<ID>IN_0</ID>236 </input>
<output>
<ID>OUT_0</ID>245 </output>
<input>
<ID>clock</ID>264 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>302</ID>
<type>AE_DFF_LOW</type>
<position>-67,183</position>
<input>
<ID>IN_0</ID>239 </input>
<output>
<ID>OUT_0</ID>248 </output>
<input>
<ID>clock</ID>264 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>304</ID>
<type>EE_VDD</type>
<position>-67.5,260.5</position>
<output>
<ID>OUT_0</ID>240 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>305</ID>
<type>AE_DFF_LOW</type>
<position>-59,237</position>
<input>
<ID>IN_0</ID>242 </input>
<output>
<ID>OUT_0</ID>367 </output>
<input>
<ID>clock</ID>249 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>306</ID>
<type>AE_DFF_LOW</type>
<position>-59,228</position>
<input>
<ID>IN_0</ID>243 </input>
<output>
<ID>OUT_0</ID>368 </output>
<input>
<ID>clock</ID>249 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>307</ID>
<type>AE_DFF_LOW</type>
<position>-59,246</position>
<input>
<ID>IN_0</ID>241 </input>
<output>
<ID>OUT_0</ID>366 </output>
<input>
<ID>clock</ID>249 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>308</ID>
<type>AE_DFF_LOW</type>
<position>-59,219</position>
<input>
<ID>IN_0</ID>244 </input>
<output>
<ID>OUT_0</ID>369 </output>
<input>
<ID>clock</ID>249 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>309</ID>
<type>AE_DFF_LOW</type>
<position>-59,201</position>
<input>
<ID>IN_0</ID>246 </input>
<output>
<ID>OUT_0</ID>371 </output>
<input>
<ID>clock</ID>249 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>310</ID>
<type>AE_DFF_LOW</type>
<position>-59,192</position>
<input>
<ID>IN_0</ID>247 </input>
<output>
<ID>OUT_0</ID>372 </output>
<input>
<ID>clock</ID>249 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>311</ID>
<type>AE_DFF_LOW</type>
<position>-59,210</position>
<input>
<ID>IN_0</ID>245 </input>
<output>
<ID>OUT_0</ID>370 </output>
<input>
<ID>clock</ID>249 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>312</ID>
<type>AE_DFF_LOW</type>
<position>-59,183</position>
<input>
<ID>IN_0</ID>248 </input>
<output>
<ID>OUT_0</ID>373 </output>
<input>
<ID>clock</ID>249 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>314</ID>
<type>DA_FROM</type>
<position>-66,178</position>
<input>
<ID>IN_0</ID>249 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>315</ID>
<type>DA_FROM</type>
<position>-74,178</position>
<input>
<ID>IN_0</ID>264 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID nclk</lparam></gate>
<gate>
<ID>319</ID>
<type>HA_JUNC_2</type>
<position>-49.5,248</position>
<input>
<ID>N_in0</ID>366 </input>
<input>
<ID>N_in1</ID>15 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>320</ID>
<type>HA_JUNC_2</type>
<position>-49.5,239</position>
<input>
<ID>N_in0</ID>367 </input>
<input>
<ID>N_in1</ID>16 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>321</ID>
<type>HA_JUNC_2</type>
<position>-49.5,230</position>
<input>
<ID>N_in0</ID>368 </input>
<input>
<ID>N_in1</ID>17 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>322</ID>
<type>HA_JUNC_2</type>
<position>-49.5,221</position>
<input>
<ID>N_in0</ID>369 </input>
<input>
<ID>N_in1</ID>18 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>323</ID>
<type>HA_JUNC_2</type>
<position>-49.5,212</position>
<input>
<ID>N_in0</ID>370 </input>
<input>
<ID>N_in1</ID>19 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>324</ID>
<type>HA_JUNC_2</type>
<position>-49.5,203</position>
<input>
<ID>N_in0</ID>371 </input>
<input>
<ID>N_in1</ID>20 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>325</ID>
<type>HA_JUNC_2</type>
<position>-49.5,194</position>
<input>
<ID>N_in0</ID>372 </input>
<input>
<ID>N_in1</ID>21 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>326</ID>
<type>HA_JUNC_2</type>
<position>-49.5,185</position>
<input>
<ID>N_in0</ID>373 </input>
<input>
<ID>N_in1</ID>22 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>345</ID>
<type>HA_JUNC_2</type>
<position>-32,212.5</position>
<input>
<ID>N_in0</ID>56 </input>
<input>
<ID>N_in1</ID>63 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>346</ID>
<type>DA_AND8</type>
<position>5,207</position>
<input>
<ID>IN_0</ID>72 </input>
<input>
<ID>IN_1</ID>73 </input>
<input>
<ID>IN_2</ID>74 </input>
<input>
<ID>IN_3</ID>75 </input>
<input>
<ID>IN_4</ID>76 </input>
<input>
<ID>IN_5</ID>79 </input>
<input>
<ID>IN_6</ID>78 </input>
<input>
<ID>IN_7</ID>77 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>372</ID>
<type>AE_OR2</type>
<position>-65.5,266</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>358 </input>
<output>
<ID>OUT</ID>334 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>373</ID>
<type>AE_OR2</type>
<position>-69.5,266</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>359 </input>
<output>
<ID>OUT</ID>335 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>374</ID>
<type>AE_OR2</type>
<position>-73.5,266</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>360 </input>
<output>
<ID>OUT</ID>336 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>375</ID>
<type>AE_OR2</type>
<position>-77.5,266</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>361 </input>
<output>
<ID>OUT</ID>337 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>377</ID>
<type>AE_OR2</type>
<position>-82.5,266</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>362 </input>
<output>
<ID>OUT</ID>333 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>378</ID>
<type>AE_OR2</type>
<position>-86.5,266</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>363 </input>
<output>
<ID>OUT</ID>338 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>379</ID>
<type>AE_OR2</type>
<position>-90.5,266</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>365 </input>
<output>
<ID>OUT</ID>339 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>380</ID>
<type>AE_OR2</type>
<position>-94.5,266</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>364 </input>
<output>
<ID>OUT</ID>340 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>382</ID>
<type>AA_AND2</type>
<position>-95.5,277</position>
<input>
<ID>IN_0</ID>375 </input>
<input>
<ID>IN_1</ID>373 </input>
<output>
<ID>OUT</ID>364 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>383</ID>
<type>AA_AND2</type>
<position>-91.5,277</position>
<input>
<ID>IN_0</ID>375 </input>
<input>
<ID>IN_1</ID>372 </input>
<output>
<ID>OUT</ID>365 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>384</ID>
<type>AA_AND2</type>
<position>-87.5,277</position>
<input>
<ID>IN_0</ID>375 </input>
<input>
<ID>IN_1</ID>371 </input>
<output>
<ID>OUT</ID>363 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>385</ID>
<type>AA_AND2</type>
<position>-83.5,277</position>
<input>
<ID>IN_0</ID>375 </input>
<input>
<ID>IN_1</ID>370 </input>
<output>
<ID>OUT</ID>362 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>386</ID>
<type>AA_AND2</type>
<position>-78.5,277</position>
<input>
<ID>IN_0</ID>375 </input>
<input>
<ID>IN_1</ID>369 </input>
<output>
<ID>OUT</ID>361 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>387</ID>
<type>AA_AND2</type>
<position>-74.5,277</position>
<input>
<ID>IN_0</ID>375 </input>
<input>
<ID>IN_1</ID>368 </input>
<output>
<ID>OUT</ID>360 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>388</ID>
<type>AA_AND2</type>
<position>-70.5,277</position>
<input>
<ID>IN_0</ID>375 </input>
<input>
<ID>IN_1</ID>367 </input>
<output>
<ID>OUT</ID>359 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-64.5,269,-64.5,269.5</points>
<connection>
<GID>372</GID>
<name>IN_0</name></connection>
<intersection>269.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-31,244,-31,269.5</points>
<connection>
<GID>428</GID>
<name>N_in1</name></connection>
<intersection>269.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-64.5,269.5,-31,269.5</points>
<intersection>-64.5 0</intersection>
<intersection>-31 1</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-68.5,269,-68.5,270</points>
<connection>
<GID>373</GID>
<name>IN_0</name></connection>
<intersection>270 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-30.5,245,-30.5,270</points>
<intersection>245 3</intersection>
<intersection>270 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-68.5,270,-30.5,270</points>
<intersection>-68.5 0</intersection>
<intersection>-30.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-30.5,245,-22.5,245</points>
<intersection>-30.5 1</intersection>
<intersection>-22.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-22.5,244.5,-22.5,245</points>
<connection>
<GID>434</GID>
<name>N_in1</name></connection>
<intersection>245 3</intersection></vsegment></shape></wire>
<wire>
<ID>391</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,306,30,306.5</points>
<connection>
<GID>420</GID>
<name>N_in1</name></connection>
<intersection>306.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>29,306.5,30,306.5</points>
<connection>
<GID>408</GID>
<name>IN_0</name></connection>
<intersection>30 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-72.5,269,-72.5,270.5</points>
<connection>
<GID>374</GID>
<name>IN_0</name></connection>
<intersection>270.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-30,245.5,-30,270.5</points>
<intersection>245.5 3</intersection>
<intersection>270.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-72.5,270.5,-30,270.5</points>
<intersection>-72.5 0</intersection>
<intersection>-30 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-30,245.5,-14,245.5</points>
<intersection>-30 1</intersection>
<intersection>-14 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-14,245,-14,245.5</points>
<connection>
<GID>439</GID>
<name>N_in1</name></connection>
<intersection>245.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>392</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,306,34,306.5</points>
<connection>
<GID>421</GID>
<name>N_in1</name></connection>
<intersection>306.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>34,306.5,35,306.5</points>
<connection>
<GID>409</GID>
<name>IN_1</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-76.5,269,-76.5,271</points>
<connection>
<GID>375</GID>
<name>IN_0</name></connection>
<intersection>271 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-29.5,246,-29.5,271</points>
<intersection>246 3</intersection>
<intersection>271 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-76.5,271,-29.5,271</points>
<intersection>-76.5 0</intersection>
<intersection>-29.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-29.5,246,-5.5,246</points>
<intersection>-29.5 1</intersection>
<intersection>-5.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-5.5,245.5,-5.5,246</points>
<connection>
<GID>444</GID>
<name>N_in1</name></connection>
<intersection>246 3</intersection></vsegment></shape></wire>
<wire>
<ID>393</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,303.5,30,304</points>
<connection>
<GID>420</GID>
<name>N_in0</name></connection>
<connection>
<GID>423</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-81.5,269,-81.5,271.5</points>
<connection>
<GID>377</GID>
<name>IN_0</name></connection>
<intersection>271.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-29,246.5,-29,271.5</points>
<intersection>246.5 3</intersection>
<intersection>271.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-81.5,271.5,-29,271.5</points>
<intersection>-81.5 0</intersection>
<intersection>-29 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-29,246.5,3,246.5</points>
<intersection>-29 1</intersection>
<intersection>3 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>3,246,3,246.5</points>
<connection>
<GID>449</GID>
<name>N_in1</name></connection>
<intersection>246.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>394</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,303.5,34,304</points>
<connection>
<GID>421</GID>
<name>N_in0</name></connection>
<connection>
<GID>425</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-85.5,269,-85.5,272</points>
<connection>
<GID>378</GID>
<name>IN_0</name></connection>
<intersection>272 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-28.5,247,-28.5,272</points>
<intersection>247 3</intersection>
<intersection>272 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-85.5,272,-28.5,272</points>
<intersection>-85.5 0</intersection>
<intersection>-28.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-28.5,247,11.5,247</points>
<intersection>-28.5 1</intersection>
<intersection>11.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>11.5,246.5,11.5,247</points>
<connection>
<GID>454</GID>
<name>N_in1</name></connection>
<intersection>247 3</intersection></vsegment></shape></wire>
<wire>
<ID>395</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,235.5,-29,241.5</points>
<intersection>235.5 3</intersection>
<intersection>241.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-31,241.5,-29,241.5</points>
<connection>
<GID>426</GID>
<name>OUT</name></connection>
<intersection>-31 31</intersection>
<intersection>-29 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-29,235.5,-28,235.5</points>
<connection>
<GID>427</GID>
<name>IN_0</name></connection>
<intersection>-29 0</intersection></hsegment>
<vsegment>
<ID>31</ID>
<points>-31,241.5,-31,242</points>
<connection>
<GID>428</GID>
<name>N_in0</name></connection>
<intersection>241.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-89.5,269,-89.5,272.5</points>
<connection>
<GID>379</GID>
<name>IN_0</name></connection>
<intersection>272.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-28,247.5,-28,272.5</points>
<intersection>247.5 3</intersection>
<intersection>272.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-89.5,272.5,-28,272.5</points>
<intersection>-89.5 0</intersection>
<intersection>-28 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-28,247.5,20,247.5</points>
<intersection>-28 1</intersection>
<intersection>20 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>20,247,20,247.5</points>
<connection>
<GID>459</GID>
<name>N_in1</name></connection>
<intersection>247.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>396</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,235.5,-29,241.5</points>
<intersection>235.5 5</intersection>
<intersection>241.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-29,241.5,-27,241.5</points>
<connection>
<GID>427</GID>
<name>OUT</name></connection>
<intersection>-29 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-30,235.5,-29,235.5</points>
<connection>
<GID>426</GID>
<name>IN_1</name></connection>
<intersection>-29 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-93.5,269,-93.5,273</points>
<connection>
<GID>380</GID>
<name>IN_0</name></connection>
<intersection>273 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-27.5,248,-27.5,273</points>
<intersection>248 3</intersection>
<intersection>273 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-93.5,273,-27.5,273</points>
<intersection>-93.5 0</intersection>
<intersection>-27.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-27.5,248,28.5,248</points>
<intersection>-27.5 1</intersection>
<intersection>28.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>28.5,247.5,28.5,248</points>
<connection>
<GID>464</GID>
<name>N_in1</name></connection>
<intersection>248 3</intersection></vsegment></shape></wire>
<wire>
<ID>397</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>-32,235.5,-31,235.5</points>
<connection>
<GID>426</GID>
<name>IN_0</name></connection>
<intersection>-31 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-31,235,-31,235.5</points>
<connection>
<GID>430</GID>
<name>N_in1</name></connection>
<intersection>235.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10.5,213.5,10.5,221.5</points>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection>
<intersection>214 56</intersection>
<intersection>214.5 53</intersection>
<intersection>221.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-26,221.5,36,221.5</points>
<intersection>-26 51</intersection>
<intersection>-17.5 4</intersection>
<intersection>-9 11</intersection>
<intersection>-0.5 13</intersection>
<intersection>8 15</intersection>
<intersection>10.5 0</intersection>
<intersection>16.5 17</intersection>
<intersection>25 19</intersection>
<intersection>33.5 21</intersection>
<intersection>36 37</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-17.5,221.5,-17.5,227</points>
<connection>
<GID>469</GID>
<name>IN_1</name></connection>
<intersection>221.5 3</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>-9,221.5,-9,227.5</points>
<connection>
<GID>470</GID>
<name>IN_1</name></connection>
<intersection>221.5 3</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>-0.5,221.5,-0.5,228</points>
<connection>
<GID>471</GID>
<name>IN_1</name></connection>
<intersection>221.5 3</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>8,221.5,8,228.5</points>
<connection>
<GID>472</GID>
<name>IN_1</name></connection>
<intersection>221.5 3</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>16.5,221.5,16.5,229</points>
<connection>
<GID>473</GID>
<name>IN_1</name></connection>
<intersection>221.5 3</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>25,221.5,25,229.5</points>
<connection>
<GID>474</GID>
<name>IN_1</name></connection>
<intersection>221.5 3</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>33.5,221.5,33.5,230</points>
<connection>
<GID>475</GID>
<name>IN_1</name></connection>
<intersection>221.5 3</intersection></vsegment>
<vsegment>
<ID>37</ID>
<points>36,221.5,36,222</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>221.5 3</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>-26,221.5,-26,226.5</points>
<connection>
<GID>468</GID>
<name>IN_1</name></connection>
<intersection>221.5 3</intersection></vsegment>
<hsegment>
<ID>53</ID>
<points>10.5,214.5,35,214.5</points>
<intersection>10.5 0</intersection>
<intersection>35 60</intersection></hsegment>
<hsegment>
<ID>56</ID>
<points>10.5,214,17,214</points>
<intersection>10.5 0</intersection>
<intersection>17 58</intersection></hsegment>
<vsegment>
<ID>58</ID>
<points>17,207.5,17,214</points>
<intersection>207.5 62</intersection>
<intersection>214 56</intersection></vsegment>
<vsegment>
<ID>60</ID>
<points>35,204,35,214.5</points>
<intersection>204 61</intersection>
<intersection>214.5 53</intersection></vsegment>
<hsegment>
<ID>61</ID>
<points>7,204,35,204</points>
<intersection>7 63</intersection>
<intersection>35 60</intersection></hsegment>
<hsegment>
<ID>62</ID>
<points>17,207.5,19.5,207.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>17 58</intersection></hsegment>
<vsegment>
<ID>63</ID>
<points>7,201,7,204</points>
<intersection>201 64</intersection>
<intersection>204 61</intersection></vsegment>
<hsegment>
<ID>64</ID>
<points>2,201,7,201</points>
<connection>
<GID>55</GID>
<name>IN_2</name></connection>
<intersection>7 63</intersection></hsegment></shape></wire>
<wire>
<ID>398</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>-27,235.5,-26,235.5</points>
<connection>
<GID>427</GID>
<name>IN_1</name></connection>
<intersection>-27 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-27,235,-27,235.5</points>
<connection>
<GID>431</GID>
<name>N_in1</name></connection>
<intersection>235.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,208,26,218</points>
<intersection>208 19</intersection>
<intersection>214 27</intersection>
<intersection>215 23</intersection>
<intersection>218 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>26,218,38,218</points>
<intersection>26 0</intersection>
<intersection>38 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>38,218,38,222</points>
<connection>
<GID>5</GID>
<name>IN_1</name></connection>
<intersection>218 2</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>26,208,28.5,208</points>
<intersection>26 0</intersection>
<intersection>28.5 22</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>28.5,207.5,28.5,208</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>208 19</intersection></vsegment>
<hsegment>
<ID>23</ID>
<points>26,215,35.5,215</points>
<intersection>26 0</intersection>
<intersection>35.5 25</intersection></hsegment>
<vsegment>
<ID>25</ID>
<points>35.5,203.5,35.5,215</points>
<intersection>203.5 26</intersection>
<intersection>215 23</intersection></vsegment>
<hsegment>
<ID>26</ID>
<points>7.5,203.5,35.5,203.5</points>
<intersection>7.5 29</intersection>
<intersection>35.5 25</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>19.5,214,26,214</points>
<intersection>19.5 28</intersection>
<intersection>26 0</intersection></hsegment>
<vsegment>
<ID>28</ID>
<points>19.5,213.5,19.5,214</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>214 27</intersection></vsegment>
<vsegment>
<ID>29</ID>
<points>7.5,199,7.5,203.5</points>
<intersection>199 30</intersection>
<intersection>203.5 26</intersection></vsegment>
<hsegment>
<ID>30</ID>
<points>2,199,7.5,199</points>
<connection>
<GID>55</GID>
<name>IN_1</name></connection>
<intersection>7.5 29</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,228,37,228.5</points>
<connection>
<GID>5</GID>
<name>OUT</name></connection>
<connection>
<GID>393</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-31,220.5,-31,233</points>
<connection>
<GID>430</GID>
<name>N_in0</name></connection>
<intersection>220.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-31,220.5,28.5,220.5</points>
<intersection>-31 0</intersection>
<intersection>-22.5 4</intersection>
<intersection>-14 6</intersection>
<intersection>-5.5 8</intersection>
<intersection>3.5 10</intersection>
<intersection>11.5 12</intersection>
<intersection>20 14</intersection>
<intersection>28.5 16</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-22.5,220.5,-22.5,233.5</points>
<connection>
<GID>435</GID>
<name>N_in0</name></connection>
<intersection>220.5 2</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-14,220.5,-14,234</points>
<connection>
<GID>440</GID>
<name>N_in0</name></connection>
<intersection>220.5 2</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>-5.5,220.5,-5.5,234.5</points>
<connection>
<GID>445</GID>
<name>N_in0</name></connection>
<intersection>220.5 2</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>3.5,220.5,3.5,235</points>
<intersection>220.5 2</intersection>
<intersection>235 27</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>11.5,220.5,11.5,235.5</points>
<connection>
<GID>455</GID>
<name>N_in0</name></connection>
<intersection>220.5 2</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>20,220.5,20,236</points>
<connection>
<GID>460</GID>
<name>N_in0</name></connection>
<intersection>220.5 2</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>28.5,213.5,28.5,236.5</points>
<connection>
<GID>465</GID>
<name>N_in0</name></connection>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>215.5 33</intersection>
<intersection>220.5 2</intersection></vsegment>
<hsegment>
<ID>27</ID>
<points>3,235,3.5,235</points>
<connection>
<GID>450</GID>
<name>N_in0</name></connection>
<intersection>3.5 10</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>28.5,215.5,36,215.5</points>
<intersection>28.5 16</intersection>
<intersection>36 34</intersection></hsegment>
<vsegment>
<ID>34</ID>
<points>36,203,36,215.5</points>
<intersection>203 35</intersection>
<intersection>215.5 33</intersection></vsegment>
<hsegment>
<ID>35</ID>
<points>8,203,36,203</points>
<intersection>8 36</intersection>
<intersection>36 34</intersection></hsegment>
<vsegment>
<ID>36</ID>
<points>8,197,8,203</points>
<intersection>197 37</intersection>
<intersection>203 35</intersection></vsegment>
<hsegment>
<ID>37</ID>
<points>2,197,8,197</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>8 36</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>13.5,205.5,13.5,207.5</points>
<connection>
<GID>1</GID>
<name>clock</name></connection>
<intersection>205.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>13.5,205.5,31.5,205.5</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>13.5 1</intersection>
<intersection>22.5 30</intersection>
<intersection>31.5 31</intersection></hsegment>
<vsegment>
<ID>30</ID>
<points>22.5,205.5,22.5,207.5</points>
<connection>
<GID>2</GID>
<name>clock</name></connection>
<intersection>205.5 2</intersection></vsegment>
<vsegment>
<ID>31</ID>
<points>31.5,205.5,31.5,207.5</points>
<connection>
<GID>3</GID>
<name>clock</name></connection>
<intersection>205.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>8,207,10.5,207</points>
<connection>
<GID>346</GID>
<name>OUT</name></connection>
<intersection>10.5 20</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>10.5,207,10.5,207.5</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<intersection>207 3</intersection></vsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-48.5,248,-44.5,248</points>
<connection>
<GID>319</GID>
<name>N_in1</name></connection>
<connection>
<GID>11</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-48,239,-48,249</points>
<intersection>239 2</intersection>
<intersection>249 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-48,249,-44.5,249</points>
<connection>
<GID>12</GID>
<name>N_in0</name></connection>
<intersection>-48 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-48.5,239,-48,239</points>
<connection>
<GID>320</GID>
<name>N_in1</name></connection>
<intersection>-48 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-47.5,230,-47.5,250</points>
<intersection>230 2</intersection>
<intersection>250 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-47.5,250,-44.5,250</points>
<connection>
<GID>13</GID>
<name>N_in0</name></connection>
<intersection>-47.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-48.5,230,-47.5,230</points>
<connection>
<GID>321</GID>
<name>N_in1</name></connection>
<intersection>-47.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-47,221,-47,251</points>
<intersection>221 2</intersection>
<intersection>251 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-47,251,-44.5,251</points>
<connection>
<GID>14</GID>
<name>N_in0</name></connection>
<intersection>-47 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-48.5,221,-47,221</points>
<connection>
<GID>322</GID>
<name>N_in1</name></connection>
<intersection>-47 0</intersection></hsegment></shape></wire>
<wire>
<ID>407</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-20.5,236,-20.5,242</points>
<intersection>236 3</intersection>
<intersection>242 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-22.5,242,-20.5,242</points>
<connection>
<GID>432</GID>
<name>OUT</name></connection>
<intersection>-22.5 32</intersection>
<intersection>-20.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-20.5,236,-19.5,236</points>
<connection>
<GID>433</GID>
<name>IN_0</name></connection>
<intersection>-20.5 0</intersection></hsegment>
<vsegment>
<ID>32</ID>
<points>-22.5,242,-22.5,242.5</points>
<connection>
<GID>434</GID>
<name>N_in0</name></connection>
<intersection>242 2</intersection></vsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46.5,212,-46.5,252</points>
<intersection>212 1</intersection>
<intersection>252 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-48.5,212,-46.5,212</points>
<connection>
<GID>323</GID>
<name>N_in1</name></connection>
<intersection>-46.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-46.5,252,-44.5,252</points>
<connection>
<GID>15</GID>
<name>N_in0</name></connection>
<intersection>-46.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>408</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-20.5,236,-20.5,242</points>
<intersection>236 5</intersection>
<intersection>242 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-20.5,242,-18.5,242</points>
<connection>
<GID>433</GID>
<name>OUT</name></connection>
<intersection>-20.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-21.5,236,-20.5,236</points>
<connection>
<GID>432</GID>
<name>IN_1</name></connection>
<intersection>-20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46,203,-46,253</points>
<intersection>203 1</intersection>
<intersection>253 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-48.5,203,-46,203</points>
<connection>
<GID>324</GID>
<name>N_in1</name></connection>
<intersection>-46 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-46,253,-44.5,253</points>
<connection>
<GID>16</GID>
<name>N_in0</name></connection>
<intersection>-46 0</intersection></hsegment></shape></wire>
<wire>
<ID>409</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>-23.5,236,-22.5,236</points>
<connection>
<GID>432</GID>
<name>IN_0</name></connection>
<intersection>-22.5 16</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>-22.5,235.5,-22.5,236</points>
<connection>
<GID>435</GID>
<name>N_in1</name></connection>
<intersection>236 4</intersection></vsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-45.5,194,-45.5,254</points>
<intersection>194 1</intersection>
<intersection>254 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-48.5,194,-45.5,194</points>
<connection>
<GID>325</GID>
<name>N_in1</name></connection>
<intersection>-45.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-45.5,254,-44.5,254</points>
<connection>
<GID>17</GID>
<name>N_in0</name></connection>
<intersection>-45.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>410</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>-18.5,236,-17.5,236</points>
<connection>
<GID>433</GID>
<name>IN_1</name></connection>
<intersection>-18.5 16</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>-18.5,235.5,-18.5,236</points>
<connection>
<GID>436</GID>
<name>N_in1</name></connection>
<intersection>236 4</intersection></vsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-45,185,-45,255</points>
<intersection>185 1</intersection>
<intersection>255 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-48.5,185,-45,185</points>
<connection>
<GID>326</GID>
<name>N_in1</name></connection>
<intersection>-45 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-45,255,-44.5,255</points>
<connection>
<GID>18</GID>
<name>N_in0</name></connection>
<intersection>-45 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36,244.5,-36,244.5</points>
<connection>
<GID>9</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>25</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,244.5,-34,244.5</points>
<connection>
<GID>9</GID>
<name>DATA_OUT_0</name></connection>
<connection>
<GID>27</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>413</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12,236.5,-12,242.5</points>
<intersection>236.5 3</intersection>
<intersection>242.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-14,242.5,-12,242.5</points>
<connection>
<GID>437</GID>
<name>OUT</name></connection>
<intersection>-14 31</intersection>
<intersection>-12 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-12,236.5,-11,236.5</points>
<connection>
<GID>438</GID>
<name>IN_0</name></connection>
<intersection>-12 0</intersection></hsegment>
<vsegment>
<ID>31</ID>
<points>-14,242.5,-14,243</points>
<connection>
<GID>439</GID>
<name>N_in0</name></connection>
<intersection>242.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35,244.5,-35,244.5</points>
<connection>
<GID>9</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>26</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>414</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12,236.5,-12,242.5</points>
<intersection>236.5 5</intersection>
<intersection>242.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-12,242.5,-10,242.5</points>
<connection>
<GID>438</GID>
<name>OUT</name></connection>
<intersection>-12 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-13,236.5,-12,236.5</points>
<connection>
<GID>437</GID>
<name>IN_1</name></connection>
<intersection>-12 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-39,244.5,-39,244.5</points>
<connection>
<GID>9</GID>
<name>DATA_OUT_5</name></connection>
<connection>
<GID>22</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>415</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>-15,236.5,-14,236.5</points>
<connection>
<GID>437</GID>
<name>IN_0</name></connection>
<intersection>-14 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-14,236,-14,236.5</points>
<connection>
<GID>440</GID>
<name>N_in1</name></connection>
<intersection>236.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-38,244.5,-38,244.5</points>
<connection>
<GID>9</GID>
<name>DATA_OUT_4</name></connection>
<connection>
<GID>23</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>416</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>-10,236.5,-9,236.5</points>
<connection>
<GID>438</GID>
<name>IN_1</name></connection>
<intersection>-10 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-10,236,-10,236.5</points>
<connection>
<GID>441</GID>
<name>N_in1</name></connection>
<intersection>236.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37,244.5,-37,244.5</points>
<connection>
<GID>9</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>24</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42.5,249,-42.5,249</points>
<connection>
<GID>9</GID>
<name>ADDRESS_1</name></connection>
<connection>
<GID>12</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>418</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3.5,237,-3.5,243</points>
<intersection>237 3</intersection>
<intersection>243 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-5.5,243,-3.5,243</points>
<connection>
<GID>442</GID>
<name>OUT</name></connection>
<intersection>-5.5 33</intersection>
<intersection>-3.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-3.5,237,-2.5,237</points>
<connection>
<GID>443</GID>
<name>IN_0</name></connection>
<intersection>-3.5 0</intersection></hsegment>
<vsegment>
<ID>33</ID>
<points>-5.5,243,-5.5,243.5</points>
<connection>
<GID>444</GID>
<name>N_in0</name></connection>
<intersection>243 2</intersection></vsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42.5,252,-42.5,252</points>
<connection>
<GID>9</GID>
<name>ADDRESS_4</name></connection>
<connection>
<GID>15</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>419</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3.5,237,-3.5,243</points>
<intersection>237 5</intersection>
<intersection>243 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-3.5,243,-1.5,243</points>
<connection>
<GID>443</GID>
<name>OUT</name></connection>
<intersection>-3.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-4.5,237,-3.5,237</points>
<connection>
<GID>442</GID>
<name>IN_1</name></connection>
<intersection>-3.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42.5,254,-42.5,254</points>
<connection>
<GID>9</GID>
<name>ADDRESS_6</name></connection>
<connection>
<GID>17</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>420</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>-6.5,237,-5.5,237</points>
<connection>
<GID>442</GID>
<name>IN_0</name></connection>
<intersection>-5.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-5.5,236.5,-5.5,237</points>
<connection>
<GID>445</GID>
<name>N_in1</name></connection>
<intersection>237 4</intersection></vsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42.5,250,-42.5,250</points>
<connection>
<GID>9</GID>
<name>ADDRESS_2</name></connection>
<connection>
<GID>13</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>421</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>-1.5,237,-0.5,237</points>
<connection>
<GID>443</GID>
<name>IN_1</name></connection>
<intersection>-1.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-1.5,236.5,-1.5,237</points>
<connection>
<GID>446</GID>
<name>N_in1</name></connection>
<intersection>237 4</intersection></vsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42.5,255,-42.5,255</points>
<connection>
<GID>9</GID>
<name>ADDRESS_7</name></connection>
<connection>
<GID>18</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-40,244.5,-40,244.5</points>
<connection>
<GID>9</GID>
<name>DATA_OUT_6</name></connection>
<connection>
<GID>21</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>423</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,237.5,5,243.5</points>
<intersection>237.5 3</intersection>
<intersection>243.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>3,243.5,5,243.5</points>
<connection>
<GID>447</GID>
<name>OUT</name></connection>
<intersection>3 15</intersection>
<intersection>5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>5,237.5,6,237.5</points>
<connection>
<GID>448</GID>
<name>IN_0</name></connection>
<intersection>5 0</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>3,243.5,3,244</points>
<connection>
<GID>449</GID>
<name>N_in0</name></connection>
<intersection>243.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42.5,253,-42.5,253</points>
<connection>
<GID>9</GID>
<name>ADDRESS_5</name></connection>
<connection>
<GID>16</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>424</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5,237.5,5,243.5</points>
<intersection>237.5 5</intersection>
<intersection>243.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>5,243.5,7,243.5</points>
<connection>
<GID>448</GID>
<name>OUT</name></connection>
<intersection>5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>4,237.5,5,237.5</points>
<connection>
<GID>447</GID>
<name>IN_1</name></connection>
<intersection>5 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-41,244.5,-41,244.5</points>
<connection>
<GID>9</GID>
<name>DATA_OUT_7</name></connection>
<connection>
<GID>20</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>425</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>2,237.5,3,237.5</points>
<connection>
<GID>447</GID>
<name>IN_0</name></connection>
<intersection>3 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>3,237,3,237.5</points>
<connection>
<GID>450</GID>
<name>N_in1</name></connection>
<intersection>237.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42.5,251,-42.5,251</points>
<connection>
<GID>9</GID>
<name>ADDRESS_3</name></connection>
<connection>
<GID>14</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>426</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>7,237.5,8,237.5</points>
<connection>
<GID>448</GID>
<name>IN_1</name></connection>
<intersection>7 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>7,237,7,237.5</points>
<connection>
<GID>451</GID>
<name>N_in1</name></connection>
<intersection>237.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42.5,248,-42.5,248</points>
<connection>
<GID>9</GID>
<name>ADDRESS_0</name></connection>
<connection>
<GID>11</GID>
<name>N_in1</name></connection></vsegment></shape></wire>
<wire>
<ID>427</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13.5,238,13.5,244</points>
<intersection>238 3</intersection>
<intersection>244 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>11.5,244,13.5,244</points>
<connection>
<GID>452</GID>
<name>OUT</name></connection>
<intersection>11.5 22</intersection>
<intersection>13.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>13.5,238,14.5,238</points>
<connection>
<GID>453</GID>
<name>IN_0</name></connection>
<intersection>13.5 0</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>11.5,244,11.5,244.5</points>
<connection>
<GID>454</GID>
<name>N_in0</name></connection>
<intersection>244 2</intersection></vsegment></shape></wire>
<wire>
<ID>428</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13.5,238,13.5,244</points>
<intersection>238 5</intersection>
<intersection>244 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>13.5,244,15.5,244</points>
<connection>
<GID>453</GID>
<name>OUT</name></connection>
<intersection>13.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>12.5,238,13.5,238</points>
<connection>
<GID>452</GID>
<name>IN_1</name></connection>
<intersection>13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-32.5,251,-31.5,251</points>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection>
<connection>
<GID>9</GID>
<name>ENABLE_0</name></connection></hsegment></shape></wire>
<wire>
<ID>429</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>10.5,238,11.5,238</points>
<connection>
<GID>452</GID>
<name>IN_0</name></connection>
<intersection>11.5 16</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>11.5,237.5,11.5,238</points>
<connection>
<GID>455</GID>
<name>N_in1</name></connection>
<intersection>238 4</intersection></vsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-31,214.5,-19,214.5</points>
<connection>
<GID>33</GID>
<name>N_in1</name></connection>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>-30 16</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>-30,214.5,-30,219.5</points>
<intersection>214.5 1</intersection>
<intersection>219.5 17</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>-30,219.5,-28,219.5</points>
<intersection>-30 16</intersection>
<intersection>-28 18</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>-28,219.5,-28,226.5</points>
<connection>
<GID>468</GID>
<name>IN_0</name></connection>
<intersection>219.5 17</intersection></vsegment></shape></wire>
<wire>
<ID>430</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>15.5,238,16.5,238</points>
<connection>
<GID>453</GID>
<name>IN_1</name></connection>
<intersection>15.5 16</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>15.5,237.5,15.5,238</points>
<connection>
<GID>456</GID>
<name>N_in1</name></connection>
<intersection>238 4</intersection></vsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-31,210.5,-20.5,210.5</points>
<connection>
<GID>32</GID>
<name>N_in1</name></connection>
<intersection>-28 16</intersection>
<intersection>-20.5 19</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>-28,210.5,-28,218.5</points>
<intersection>210.5 1</intersection>
<intersection>218.5 17</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>-28,218.5,-11,218.5</points>
<intersection>-28 16</intersection>
<intersection>-11 18</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>-11,218.5,-11,227.5</points>
<connection>
<GID>470</GID>
<name>IN_0</name></connection>
<intersection>218.5 17</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>-20.5,206.5,-20.5,210.5</points>
<intersection>206.5 20</intersection>
<intersection>210.5 1</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>-20.5,206.5,-19,206.5</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>-20.5 19</intersection></hsegment></shape></wire>
<wire>
<ID>431</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,238.5,22,244.5</points>
<intersection>238.5 3</intersection>
<intersection>244.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>20,244.5,22,244.5</points>
<connection>
<GID>457</GID>
<name>OUT</name></connection>
<intersection>20 29</intersection>
<intersection>22 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>22,238.5,23,238.5</points>
<connection>
<GID>458</GID>
<name>IN_0</name></connection>
<intersection>22 0</intersection></hsegment>
<vsegment>
<ID>29</ID>
<points>20,244.5,20,245</points>
<connection>
<GID>459</GID>
<name>N_in0</name></connection>
<intersection>244.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-31,208.5,-21,208.5</points>
<connection>
<GID>37</GID>
<name>N_in1</name></connection>
<intersection>-27 8</intersection>
<intersection>-21 23</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-27,208.5,-27,218</points>
<intersection>208.5 1</intersection>
<intersection>218 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-27,218,-2.5,218</points>
<intersection>-27 8</intersection>
<intersection>-2.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-2.5,218,-2.5,228</points>
<connection>
<GID>471</GID>
<name>IN_0</name></connection>
<intersection>218 9</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>-21,202.5,-21,208.5</points>
<intersection>202.5 24</intersection>
<intersection>208.5 1</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>-21,202.5,-19,202.5</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>-21 23</intersection></hsegment></shape></wire>
<wire>
<ID>432</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,238.5,22,244.5</points>
<intersection>238.5 5</intersection>
<intersection>244.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>22,244.5,24,244.5</points>
<connection>
<GID>458</GID>
<name>OUT</name></connection>
<intersection>22 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>21,238.5,22,238.5</points>
<connection>
<GID>457</GID>
<name>IN_1</name></connection>
<intersection>22 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-31,206.5,-21.5,206.5</points>
<connection>
<GID>38</GID>
<name>N_in1</name></connection>
<intersection>-26 8</intersection>
<intersection>-21.5 23</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-26,206.5,-26,217.5</points>
<intersection>206.5 1</intersection>
<intersection>217.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-26,217.5,6,217.5</points>
<intersection>-26 8</intersection>
<intersection>6 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>6,217.5,6,228.5</points>
<connection>
<GID>472</GID>
<name>IN_0</name></connection>
<intersection>217.5 9</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>-21.5,197.5,-21.5,206.5</points>
<intersection>197.5 24</intersection>
<intersection>206.5 1</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>-21.5,197.5,-19,197.5</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>-21.5 23</intersection></hsegment></shape></wire>
<wire>
<ID>433</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>19,238.5,20,238.5</points>
<connection>
<GID>457</GID>
<name>IN_0</name></connection>
<intersection>20 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>20,238,20,238.5</points>
<connection>
<GID>460</GID>
<name>N_in1</name></connection>
<intersection>238.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-31,204.5,-22,204.5</points>
<connection>
<GID>39</GID>
<name>N_in1</name></connection>
<intersection>-25 12</intersection>
<intersection>-22 28</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>-25,204.5,-25,217</points>
<intersection>204.5 1</intersection>
<intersection>217 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>-25,217,14.5,217</points>
<intersection>-25 12</intersection>
<intersection>14.5 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>14.5,217,14.5,229</points>
<connection>
<GID>473</GID>
<name>IN_0</name></connection>
<intersection>217 13</intersection></vsegment>
<vsegment>
<ID>28</ID>
<points>-22,193.5,-22,204.5</points>
<intersection>193.5 29</intersection>
<intersection>204.5 1</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>-22,193.5,-19,193.5</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<intersection>-22 28</intersection></hsegment></shape></wire>
<wire>
<ID>434</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>24,238.5,25,238.5</points>
<connection>
<GID>458</GID>
<name>IN_1</name></connection>
<intersection>24 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>24,238,24,238.5</points>
<connection>
<GID>461</GID>
<name>N_in1</name></connection>
<intersection>238.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-31,202.5,-22.5,202.5</points>
<connection>
<GID>40</GID>
<name>N_in1</name></connection>
<intersection>-24 12</intersection>
<intersection>-22.5 27</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>-24,202.5,-24,216.5</points>
<intersection>202.5 1</intersection>
<intersection>216.5 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>-24,216.5,23,216.5</points>
<intersection>-24 12</intersection>
<intersection>23 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>23,216.5,23,229.5</points>
<connection>
<GID>474</GID>
<name>IN_0</name></connection>
<intersection>216.5 13</intersection></vsegment>
<vsegment>
<ID>27</ID>
<points>-22.5,189.5,-22.5,202.5</points>
<intersection>189.5 28</intersection>
<intersection>202.5 1</intersection></vsegment>
<hsegment>
<ID>28</ID>
<points>-22.5,189.5,-19,189.5</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>-22.5 27</intersection></hsegment></shape></wire>
<wire>
<ID>435</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,239.5,30.5,245</points>
<intersection>239.5 3</intersection>
<intersection>245 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>28.5,245,30.5,245</points>
<connection>
<GID>462</GID>
<name>OUT</name></connection>
<intersection>28.5 33</intersection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>30.5,239.5,31.5,239.5</points>
<intersection>30.5 0</intersection>
<intersection>31.5 26</intersection></hsegment>
<vsegment>
<ID>26</ID>
<points>31.5,239,31.5,239.5</points>
<connection>
<GID>463</GID>
<name>IN_0</name></connection>
<intersection>239.5 3</intersection></vsegment>
<vsegment>
<ID>33</ID>
<points>28.5,245,28.5,245.5</points>
<connection>
<GID>464</GID>
<name>N_in0</name></connection>
<intersection>245 2</intersection></vsegment></shape></wire>
<wire>
<ID>436</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,239,30.5,245</points>
<intersection>239 5</intersection>
<intersection>245 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>30.5,245,32.5,245</points>
<connection>
<GID>463</GID>
<name>OUT</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>29.5,239,30.5,239</points>
<connection>
<GID>462</GID>
<name>IN_1</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-31,200.5,-23,200.5</points>
<connection>
<GID>41</GID>
<name>N_in1</name></connection>
<intersection>-23 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>-23,185.5,-23,216</points>
<intersection>185.5 28</intersection>
<intersection>200.5 1</intersection>
<intersection>216 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>-23,216,31.5,216</points>
<intersection>-23 12</intersection>
<intersection>31.5 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>31.5,216,31.5,230</points>
<connection>
<GID>475</GID>
<name>IN_0</name></connection>
<intersection>216 13</intersection></vsegment>
<hsegment>
<ID>28</ID>
<points>-23,185.5,-19,185.5</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<intersection>-23 12</intersection></hsegment></shape></wire>
<wire>
<ID>437</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>27.5,239,28.5,239</points>
<connection>
<GID>462</GID>
<name>IN_0</name></connection>
<intersection>28.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>28.5,238.5,28.5,239</points>
<connection>
<GID>465</GID>
<name>N_in1</name></connection>
<intersection>239 4</intersection></vsegment></shape></wire>
<wire>
<ID>438</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>32.5,239,33.5,239</points>
<connection>
<GID>463</GID>
<name>IN_1</name></connection>
<intersection>32.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>32.5,238.5,32.5,239</points>
<connection>
<GID>466</GID>
<name>N_in1</name></connection>
<intersection>239 4</intersection></vsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,214.5,-34,242.5</points>
<connection>
<GID>27</GID>
<name>N_in0</name></connection>
<intersection>214.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34,214.5,-33,214.5</points>
<connection>
<GID>33</GID>
<name>N_in0</name></connection>
<intersection>-34 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35,212.5,-35,242.5</points>
<connection>
<GID>26</GID>
<name>N_in0</name></connection>
<intersection>212.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-35,212.5,-33,212.5</points>
<connection>
<GID>345</GID>
<name>N_in0</name></connection>
<intersection>-35 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36,210.5,-36,242.5</points>
<connection>
<GID>25</GID>
<name>N_in0</name></connection>
<intersection>210.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36,210.5,-33,210.5</points>
<connection>
<GID>32</GID>
<name>N_in0</name></connection>
<intersection>-36 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37,208.5,-37,242.5</points>
<connection>
<GID>24</GID>
<name>N_in0</name></connection>
<intersection>208.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-37,208.5,-33,208.5</points>
<connection>
<GID>37</GID>
<name>N_in0</name></connection>
<intersection>-37 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-38,206.5,-38,242.5</points>
<connection>
<GID>23</GID>
<name>N_in0</name></connection>
<intersection>206.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-38,206.5,-33,206.5</points>
<connection>
<GID>38</GID>
<name>N_in0</name></connection>
<intersection>-38 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-39,204.5,-39,242.5</points>
<connection>
<GID>22</GID>
<name>N_in0</name></connection>
<intersection>204.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-39,204.5,-33,204.5</points>
<connection>
<GID>39</GID>
<name>N_in0</name></connection>
<intersection>-39 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-40,202.5,-40,242.5</points>
<connection>
<GID>21</GID>
<name>N_in0</name></connection>
<intersection>202.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-40,202.5,-33,202.5</points>
<connection>
<GID>40</GID>
<name>N_in0</name></connection>
<intersection>-40 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-41,200.5,-41,242.5</points>
<connection>
<GID>20</GID>
<name>N_in0</name></connection>
<intersection>200.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-41,200.5,-33,200.5</points>
<connection>
<GID>41</GID>
<name>N_in0</name></connection>
<intersection>-41 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,212.5,-29,219</points>
<intersection>212.5 1</intersection>
<intersection>219 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-31,212.5,-20,212.5</points>
<connection>
<GID>345</GID>
<name>N_in1</name></connection>
<intersection>-29 0</intersection>
<intersection>-20 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-29,219,-19.5,219</points>
<intersection>-29 0</intersection>
<intersection>-19.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-19.5,219,-19.5,227</points>
<connection>
<GID>469</GID>
<name>IN_0</name></connection>
<intersection>219 2</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-20,210.5,-20,212.5</points>
<intersection>210.5 6</intersection>
<intersection>212.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-20,210.5,-19,210.5</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>-20 5</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13,213.5,-12,213.5</points>
<connection>
<GID>50</GID>
<name>OUT</name></connection>
<connection>
<GID>57</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13,201.5,-12,201.5</points>
<connection>
<GID>53</GID>
<name>OUT</name></connection>
<connection>
<GID>59</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13,205.5,-12,205.5</points>
<connection>
<GID>52</GID>
<name>OUT</name></connection>
<connection>
<GID>58</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13,196.5,-12,196.5</points>
<connection>
<GID>60</GID>
<name>OUT</name></connection>
<connection>
<GID>64</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>456</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-27,232.5,-27,233</points>
<connection>
<GID>468</GID>
<name>OUT</name></connection>
<connection>
<GID>431</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13,184.5,-12,184.5</points>
<connection>
<GID>63</GID>
<name>OUT</name></connection>
<connection>
<GID>66</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>457</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-18.5,233,-18.5,233.5</points>
<connection>
<GID>469</GID>
<name>OUT</name></connection>
<connection>
<GID>436</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13,188.5,-12,188.5</points>
<connection>
<GID>62</GID>
<name>OUT</name></connection>
<connection>
<GID>65</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>458</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-10,233.5,-10,234</points>
<connection>
<GID>470</GID>
<name>OUT</name></connection>
<connection>
<GID>441</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13,192.5,-12,192.5</points>
<connection>
<GID>61</GID>
<name>OUT</name></connection>
<connection>
<GID>67</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>459</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1.5,234,-1.5,234.5</points>
<connection>
<GID>471</GID>
<name>OUT</name></connection>
<connection>
<GID>446</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>460</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,234.5,7,235</points>
<connection>
<GID>472</GID>
<name>OUT</name></connection>
<connection>
<GID>451</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7,210.5,-7,213.5</points>
<intersection>210.5 1</intersection>
<intersection>213.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-7,210.5,2,210.5</points>
<connection>
<GID>346</GID>
<name>IN_0</name></connection>
<intersection>-7 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-8,213.5,-7,213.5</points>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection>
<intersection>-7 0</intersection></hsegment></shape></wire>
<wire>
<ID>461</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15.5,235,15.5,235.5</points>
<connection>
<GID>473</GID>
<name>OUT</name></connection>
<connection>
<GID>456</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13,209.5,2,209.5</points>
<connection>
<GID>51</GID>
<name>OUT</name></connection>
<connection>
<GID>346</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>462</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,235.5,24,236</points>
<connection>
<GID>474</GID>
<name>OUT</name></connection>
<connection>
<GID>461</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7,205.5,-7,208.5</points>
<intersection>205.5 2</intersection>
<intersection>208.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-7,208.5,2,208.5</points>
<connection>
<GID>346</GID>
<name>IN_2</name></connection>
<intersection>-7 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-8,205.5,-7,205.5</points>
<connection>
<GID>58</GID>
<name>OUT_0</name></connection>
<intersection>-7 0</intersection></hsegment></shape></wire>
<wire>
<ID>463</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,236,32.5,236.5</points>
<connection>
<GID>475</GID>
<name>OUT</name></connection>
<connection>
<GID>466</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6.5,201.5,-6.5,207.5</points>
<intersection>201.5 2</intersection>
<intersection>207.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-6.5,207.5,2,207.5</points>
<connection>
<GID>346</GID>
<name>IN_3</name></connection>
<intersection>-6.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-8,201.5,-6.5,201.5</points>
<connection>
<GID>59</GID>
<name>OUT_0</name></connection>
<intersection>-6.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6,196.5,-6,206.5</points>
<intersection>196.5 2</intersection>
<intersection>206.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-6,206.5,2,206.5</points>
<connection>
<GID>346</GID>
<name>IN_4</name></connection>
<intersection>-6 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-8,196.5,-6,196.5</points>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection>
<intersection>-6 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,184.5,-4.5,203.5</points>
<intersection>184.5 2</intersection>
<intersection>203.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,203.5,2,203.5</points>
<connection>
<GID>346</GID>
<name>IN_7</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-8,184.5,-4.5,184.5</points>
<connection>
<GID>66</GID>
<name>OUT_0</name></connection>
<intersection>-4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5,188.5,-5,204.5</points>
<intersection>188.5 2</intersection>
<intersection>204.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-5,204.5,2,204.5</points>
<connection>
<GID>346</GID>
<name>IN_6</name></connection>
<intersection>-5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-8,188.5,-5,188.5</points>
<connection>
<GID>65</GID>
<name>OUT_0</name></connection>
<intersection>-5 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5.5,192.5,-5.5,205.5</points>
<intersection>192.5 2</intersection>
<intersection>205.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-5.5,205.5,2,205.5</points>
<connection>
<GID>346</GID>
<name>IN_5</name></connection>
<intersection>-5.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-8,192.5,-5.5,192.5</points>
<connection>
<GID>67</GID>
<name>OUT_0</name></connection>
<intersection>-5.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-7,199,-4,199</points>
<connection>
<GID>55</GID>
<name>OUT</name></connection>
<connection>
<GID>69</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-19.5,183.5,-19.5,212.5</points>
<intersection>183.5 7</intersection>
<intersection>187.5 10</intersection>
<intersection>191.5 9</intersection>
<intersection>195.5 8</intersection>
<intersection>199 2</intersection>
<intersection>200.5 5</intersection>
<intersection>204.5 4</intersection>
<intersection>208.5 3</intersection>
<intersection>212.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-19.5,212.5,-19,212.5</points>
<connection>
<GID>50</GID>
<name>IN_1</name></connection>
<intersection>-19.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-19.5,199,-11,199</points>
<connection>
<GID>69</GID>
<name>OUT_0</name></connection>
<intersection>-19.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-19.5,208.5,-19,208.5</points>
<connection>
<GID>51</GID>
<name>IN_1</name></connection>
<intersection>-19.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-19.5,204.5,-19,204.5</points>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<intersection>-19.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-19.5,200.5,-19,200.5</points>
<connection>
<GID>53</GID>
<name>IN_1</name></connection>
<intersection>-19.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-19.5,183.5,-19,183.5</points>
<connection>
<GID>63</GID>
<name>IN_1</name></connection>
<intersection>-19.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-19.5,195.5,-19,195.5</points>
<connection>
<GID>60</GID>
<name>IN_1</name></connection>
<intersection>-19.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-19.5,191.5,-19,191.5</points>
<connection>
<GID>61</GID>
<name>IN_1</name></connection>
<intersection>-19.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-19.5,187.5,-19,187.5</points>
<connection>
<GID>62</GID>
<name>IN_1</name></connection>
<intersection>-19.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>32.5,151,32.5,153</points>
<intersection>151 5</intersection>
<intersection>153 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>29,153,32.5,153</points>
<connection>
<GID>185</GID>
<name>OUT_2</name></connection>
<intersection>32.5 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>32.5,151,33.5,151</points>
<connection>
<GID>179</GID>
<name>ADDRESS_2</name></connection>
<intersection>32.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>32,150,32,151</points>
<intersection>150 5</intersection>
<intersection>151 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>29,151,32,151</points>
<connection>
<GID>185</GID>
<name>OUT_1</name></connection>
<intersection>32 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>32,150,33.5,150</points>
<connection>
<GID>179</GID>
<name>ADDRESS_1</name></connection>
<intersection>32 3</intersection></hsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,152,33,155</points>
<intersection>152 5</intersection>
<intersection>155 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>29,155,33,155</points>
<connection>
<GID>185</GID>
<name>OUT_3</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>33,152,33.5,152</points>
<connection>
<GID>179</GID>
<name>ADDRESS_3</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29,149,33.5,149</points>
<connection>
<GID>179</GID>
<name>ADDRESS_0</name></connection>
<connection>
<GID>185</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>213</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,143,40,145.5</points>
<connection>
<GID>179</GID>
<name>DATA_OUT_0</name></connection>
<connection>
<GID>179</GID>
<name>DATA_IN_0</name></connection>
<intersection>143 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>35,142.5,35,143</points>
<connection>
<GID>203</GID>
<name>OUT</name></connection>
<intersection>143 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>35,143,54,143</points>
<intersection>35 1</intersection>
<intersection>40 0</intersection>
<intersection>54 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>54,142.5,54,143</points>
<connection>
<GID>214</GID>
<name>IN_1</name></connection>
<intersection>143 2</intersection></vsegment></shape></wire>
<wire>
<ID>214</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,143.5,39,145.5</points>
<connection>
<GID>179</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>179</GID>
<name>DATA_IN_1</name></connection>
<intersection>143.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>31,142.5,31,143.5</points>
<connection>
<GID>205</GID>
<name>OUT</name></connection>
<intersection>143.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>31,143.5,50,143.5</points>
<intersection>31 1</intersection>
<intersection>39 0</intersection>
<intersection>50 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>50,142.5,50,143.5</points>
<connection>
<GID>213</GID>
<name>IN_1</name></connection>
<intersection>143.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>215</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,144.5,37,145.5</points>
<connection>
<GID>179</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>179</GID>
<name>DATA_IN_3</name></connection>
<intersection>144.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>23,142.5,23,144.5</points>
<connection>
<GID>207</GID>
<name>OUT</name></connection>
<intersection>144.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>23,144.5,42,144.5</points>
<intersection>23 1</intersection>
<intersection>37 0</intersection>
<intersection>42 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>42,142.5,42,144.5</points>
<connection>
<GID>211</GID>
<name>IN_1</name></connection>
<intersection>144.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>216</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,144,38,145.5</points>
<connection>
<GID>179</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>179</GID>
<name>DATA_IN_2</name></connection>
<intersection>144 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>27,142.5,27,144</points>
<connection>
<GID>206</GID>
<name>OUT</name></connection>
<intersection>144 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>27,144,46,144</points>
<intersection>27 1</intersection>
<intersection>38 0</intersection>
<intersection>46 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>46,142.5,46,144</points>
<connection>
<GID>212</GID>
<name>IN_1</name></connection>
<intersection>144 2</intersection></vsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43.5,150,56,150</points>
<connection>
<GID>179</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>216</GID>
<name>OUT_0</name></connection>
<intersection>44 10</intersection>
<intersection>48 11</intersection>
<intersection>52 9</intersection>
<intersection>56 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>56,142.5,56,150</points>
<connection>
<GID>214</GID>
<name>IN_0</name></connection>
<intersection>150 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>52,142.5,52,150</points>
<connection>
<GID>213</GID>
<name>IN_0</name></connection>
<intersection>150 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>44,142.5,44,150</points>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<intersection>150 1</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>48,142.5,48,150</points>
<connection>
<GID>212</GID>
<name>IN_0</name></connection>
<intersection>150 1</intersection></vsegment></shape></wire>
<wire>
<ID>219</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,152,44.5,156.5</points>
<intersection>152 1</intersection>
<intersection>156.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,152,44.5,152</points>
<connection>
<GID>179</GID>
<name>write_clock</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>42.5,156.5,44.5,156.5</points>
<connection>
<GID>218</GID>
<name>CLK</name></connection>
<intersection>44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,133.5,51,136.5</points>
<connection>
<GID>213</GID>
<name>OUT</name></connection>
<intersection>133.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51,133.5,57,133.5</points>
<connection>
<GID>183</GID>
<name>IN_1</name></connection>
<intersection>51 0</intersection></hsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,132.5,55,136.5</points>
<connection>
<GID>214</GID>
<name>OUT</name></connection>
<intersection>132.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55,132.5,57,132.5</points>
<connection>
<GID>183</GID>
<name>IN_0</name></connection>
<intersection>55 0</intersection></hsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,134.5,47,136.5</points>
<connection>
<GID>212</GID>
<name>OUT</name></connection>
<intersection>134.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,134.5,57,134.5</points>
<connection>
<GID>183</GID>
<name>IN_2</name></connection>
<intersection>47 0</intersection></hsegment></shape></wire>
<wire>
<ID>226</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,135.5,43,136.5</points>
<connection>
<GID>211</GID>
<name>OUT</name></connection>
<intersection>135.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43,135.5,57,135.5</points>
<connection>
<GID>183</GID>
<name>IN_3</name></connection>
<intersection>43 0</intersection></hsegment></shape></wire>
<wire>
<ID>227</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19,159.5,52.5,159.5</points>
<intersection>19 4</intersection>
<intersection>52.5 6</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>19,135.5,19,159.5</points>
<intersection>135.5 10</intersection>
<intersection>159.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>52.5,151,52.5,159.5</points>
<connection>
<GID>220</GID>
<name>OUT_0</name></connection>
<intersection>151 11</intersection>
<intersection>159.5 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>19,135.5,34,135.5</points>
<intersection>19 4</intersection>
<intersection>22 12</intersection>
<intersection>26 14</intersection>
<intersection>30 16</intersection>
<intersection>34 18</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>43.5,151,52.5,151</points>
<connection>
<GID>179</GID>
<name>write_enable</name></connection>
<intersection>52.5 6</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>22,135.5,22,136.5</points>
<connection>
<GID>207</GID>
<name>IN_0</name></connection>
<intersection>135.5 10</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>26,135.5,26,136.5</points>
<connection>
<GID>206</GID>
<name>IN_0</name></connection>
<intersection>135.5 10</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>30,135.5,30,136.5</points>
<connection>
<GID>205</GID>
<name>IN_0</name></connection>
<intersection>135.5 10</intersection></vsegment>
<vsegment>
<ID>18</ID>
<points>34,135.5,34,136.5</points>
<connection>
<GID>203</GID>
<name>IN_0</name></connection>
<intersection>135.5 10</intersection></vsegment></shape></wire>
<wire>
<ID>228</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,132.5,24,136.5</points>
<connection>
<GID>207</GID>
<name>IN_1</name></connection>
<intersection>132.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15.5,132.5,24,132.5</points>
<connection>
<GID>201</GID>
<name>OUT_3</name></connection>
<intersection>24 0</intersection></hsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-81.5,256,-80.5,256</points>
<connection>
<GID>296</GID>
<name>carry_out</name></connection>
<connection>
<GID>298</GID>
<name>carry_in</name></connection></hsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-71,248,-71,251</points>
<connection>
<GID>296</GID>
<name>OUT_0</name></connection>
<intersection>248 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-71,248,-70,248</points>
<connection>
<GID>293</GID>
<name>IN_0</name></connection>
<intersection>-71 0</intersection></hsegment></shape></wire>
<wire>
<ID>231</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-72,239,-72,251</points>
<connection>
<GID>296</GID>
<name>OUT_1</name></connection>
<intersection>239 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-72,239,-70,239</points>
<connection>
<GID>290</GID>
<name>IN_0</name></connection>
<intersection>-72 0</intersection></hsegment></shape></wire>
<wire>
<ID>232</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,130.5,28,136.5</points>
<connection>
<GID>206</GID>
<name>IN_1</name></connection>
<intersection>130.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15.5,130.5,28,130.5</points>
<connection>
<GID>201</GID>
<name>OUT_2</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>233</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,128.5,32,136.5</points>
<connection>
<GID>205</GID>
<name>IN_1</name></connection>
<intersection>128.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15.5,128.5,32,128.5</points>
<connection>
<GID>201</GID>
<name>OUT_1</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>234</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-73,230,-73,251</points>
<connection>
<GID>296</GID>
<name>OUT_2</name></connection>
<intersection>230 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-73,230,-70,230</points>
<connection>
<GID>291</GID>
<name>IN_0</name></connection>
<intersection>-73 0</intersection></hsegment></shape></wire>
<wire>
<ID>235</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-74,221,-74,251</points>
<connection>
<GID>296</GID>
<name>OUT_3</name></connection>
<intersection>221 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-74,221,-70,221</points>
<connection>
<GID>294</GID>
<name>IN_0</name></connection>
<intersection>-74 0</intersection></hsegment></shape></wire>
<wire>
<ID>236</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-75,212,-75,250</points>
<intersection>212 1</intersection>
<intersection>250 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-75,212,-70,212</points>
<connection>
<GID>301</GID>
<name>IN_0</name></connection>
<intersection>-75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-88,250,-75,250</points>
<intersection>-88 3</intersection>
<intersection>-75 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-88,250,-88,251</points>
<connection>
<GID>298</GID>
<name>OUT_0</name></connection>
<intersection>250 2</intersection></vsegment></shape></wire>
<wire>
<ID>237</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-76,203,-76,249</points>
<intersection>203 1</intersection>
<intersection>249 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-76,203,-70,203</points>
<connection>
<GID>299</GID>
<name>IN_0</name></connection>
<intersection>-76 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-89,249,-76,249</points>
<intersection>-89 3</intersection>
<intersection>-76 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-89,249,-89,251</points>
<connection>
<GID>298</GID>
<name>OUT_1</name></connection>
<intersection>249 2</intersection></vsegment></shape></wire>
<wire>
<ID>238</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-77,194,-77,248</points>
<intersection>194 1</intersection>
<intersection>248 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-77,194,-70,194</points>
<connection>
<GID>300</GID>
<name>IN_0</name></connection>
<intersection>-77 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-90,248,-77,248</points>
<intersection>-90 3</intersection>
<intersection>-77 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-90,248,-90,251</points>
<connection>
<GID>298</GID>
<name>OUT_2</name></connection>
<intersection>248 2</intersection></vsegment></shape></wire>
<wire>
<ID>239</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-78,185,-78,247</points>
<intersection>185 1</intersection>
<intersection>247 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-78,185,-70,185</points>
<connection>
<GID>302</GID>
<name>IN_0</name></connection>
<intersection>-78 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-91,247,-78,247</points>
<intersection>-91 3</intersection>
<intersection>-78 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-91,247,-91,251</points>
<connection>
<GID>298</GID>
<name>OUT_3</name></connection>
<intersection>247 2</intersection></vsegment></shape></wire>
<wire>
<ID>240</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-67.5,259,-67.5,259.5</points>
<connection>
<GID>296</GID>
<name>IN_B_0</name></connection>
<connection>
<GID>304</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>241</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-64,248,-62,248</points>
<connection>
<GID>307</GID>
<name>IN_0</name></connection>
<connection>
<GID>293</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>242</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-64,239,-62,239</points>
<connection>
<GID>305</GID>
<name>IN_0</name></connection>
<connection>
<GID>290</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>243</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-64,230,-62,230</points>
<connection>
<GID>291</GID>
<name>OUT_0</name></connection>
<connection>
<GID>306</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>244</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-64,221,-62,221</points>
<connection>
<GID>308</GID>
<name>IN_0</name></connection>
<connection>
<GID>294</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>245</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-64,212,-62,212</points>
<connection>
<GID>311</GID>
<name>IN_0</name></connection>
<connection>
<GID>301</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>246</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-64,203,-62,203</points>
<connection>
<GID>309</GID>
<name>IN_0</name></connection>
<connection>
<GID>299</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>247</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-64,194,-62,194</points>
<connection>
<GID>310</GID>
<name>IN_0</name></connection>
<connection>
<GID>300</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>248</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-64,185,-62,185</points>
<connection>
<GID>312</GID>
<name>IN_0</name></connection>
<connection>
<GID>302</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>249</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63,178,-63,245</points>
<intersection>178 1</intersection>
<intersection>182 9</intersection>
<intersection>191 8</intersection>
<intersection>200 7</intersection>
<intersection>209 6</intersection>
<intersection>218 5</intersection>
<intersection>227 4</intersection>
<intersection>236 3</intersection>
<intersection>245 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-64,178,-63,178</points>
<connection>
<GID>314</GID>
<name>IN_0</name></connection>
<intersection>-63 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-63,245,-62,245</points>
<connection>
<GID>307</GID>
<name>clock</name></connection>
<intersection>-63 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-63,236,-62,236</points>
<connection>
<GID>305</GID>
<name>clock</name></connection>
<intersection>-63 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-63,227,-62,227</points>
<connection>
<GID>306</GID>
<name>clock</name></connection>
<intersection>-63 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-63,218,-62,218</points>
<connection>
<GID>308</GID>
<name>clock</name></connection>
<intersection>-63 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-63,209,-62,209</points>
<connection>
<GID>311</GID>
<name>clock</name></connection>
<intersection>-63 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-63,200,-62,200</points>
<connection>
<GID>309</GID>
<name>clock</name></connection>
<intersection>-63 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-63,191,-62,191</points>
<connection>
<GID>310</GID>
<name>clock</name></connection>
<intersection>-63 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-63,182,-62,182</points>
<connection>
<GID>312</GID>
<name>clock</name></connection>
<intersection>-63 0</intersection></hsegment></shape></wire>
<wire>
<ID>250</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,126.5,36,136.5</points>
<connection>
<GID>203</GID>
<name>IN_1</name></connection>
<intersection>126.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15.5,126.5,36,126.5</points>
<connection>
<GID>201</GID>
<name>OUT_0</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>264</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-71,178,-71,245</points>
<intersection>178 1</intersection>
<intersection>182 9</intersection>
<intersection>191 8</intersection>
<intersection>200 7</intersection>
<intersection>209 6</intersection>
<intersection>218 5</intersection>
<intersection>227 4</intersection>
<intersection>236 3</intersection>
<intersection>245 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-72,178,-71,178</points>
<connection>
<GID>315</GID>
<name>IN_0</name></connection>
<intersection>-71 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71,245,-70,245</points>
<connection>
<GID>293</GID>
<name>clock</name></connection>
<intersection>-71 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-71,236,-70,236</points>
<connection>
<GID>290</GID>
<name>clock</name></connection>
<intersection>-71 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-71,227,-70,227</points>
<connection>
<GID>291</GID>
<name>clock</name></connection>
<intersection>-71 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-71,218,-70,218</points>
<connection>
<GID>294</GID>
<name>clock</name></connection>
<intersection>-71 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-71,209,-70,209</points>
<connection>
<GID>301</GID>
<name>clock</name></connection>
<intersection>-71 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-71,200,-70,200</points>
<connection>
<GID>299</GID>
<name>clock</name></connection>
<intersection>-71 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-71,191,-70,191</points>
<connection>
<GID>300</GID>
<name>clock</name></connection>
<intersection>-71 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-71,182,-70,182</points>
<connection>
<GID>302</GID>
<name>clock</name></connection>
<intersection>-71 0</intersection></hsegment></shape></wire>
<wire>
<ID>301</ID>
<shape>
<hsegment>
<ID>11</ID>
<points>8.5,269.5,9,269.5</points>
<connection>
<GID>270</GID>
<name>OUT_0</name></connection>
<connection>
<GID>272</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>302</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4.5,267.5,4.5,269.5</points>
<connection>
<GID>270</GID>
<name>IN_0</name></connection>
<intersection>267.5 2</intersection>
<intersection>268.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3,268.5,4.5,268.5</points>
<connection>
<GID>268</GID>
<name>CLK</name></connection>
<intersection>4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>4.5,267.5,9,267.5</points>
<connection>
<GID>274</GID>
<name>IN_0</name></connection>
<intersection>4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>333</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-91.5,259,-91.5,261.5</points>
<connection>
<GID>298</GID>
<name>IN_0</name></connection>
<intersection>261.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-82.5,261.5,-82.5,263</points>
<connection>
<GID>377</GID>
<name>OUT</name></connection>
<intersection>261.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-91.5,261.5,-82.5,261.5</points>
<intersection>-91.5 0</intersection>
<intersection>-82.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>334</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-74.5,259,-74.5,261.5</points>
<connection>
<GID>296</GID>
<name>IN_0</name></connection>
<intersection>261.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-65.5,261.5,-65.5,263</points>
<connection>
<GID>372</GID>
<name>OUT</name></connection>
<intersection>261.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-74.5,261.5,-65.5,261.5</points>
<intersection>-74.5 0</intersection>
<intersection>-65.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>335</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-75.5,259,-75.5,262</points>
<connection>
<GID>296</GID>
<name>IN_1</name></connection>
<intersection>262 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-75.5,262,-69.5,262</points>
<intersection>-75.5 0</intersection>
<intersection>-69.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-69.5,262,-69.5,263</points>
<connection>
<GID>373</GID>
<name>OUT</name></connection>
<intersection>262 2</intersection></vsegment></shape></wire>
<wire>
<ID>336</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-76.5,259,-76.5,262.5</points>
<connection>
<GID>296</GID>
<name>IN_2</name></connection>
<intersection>262.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-73.5,262.5,-73.5,263</points>
<connection>
<GID>374</GID>
<name>OUT</name></connection>
<intersection>262.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-76.5,262.5,-73.5,262.5</points>
<intersection>-76.5 0</intersection>
<intersection>-73.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>337</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-77.5,259,-77.5,263</points>
<connection>
<GID>296</GID>
<name>IN_3</name></connection>
<connection>
<GID>375</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>338</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-92.5,259,-92.5,262</points>
<connection>
<GID>298</GID>
<name>IN_1</name></connection>
<intersection>262 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-86.5,262,-86.5,263</points>
<connection>
<GID>378</GID>
<name>OUT</name></connection>
<intersection>262 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-92.5,262,-86.5,262</points>
<intersection>-92.5 0</intersection>
<intersection>-86.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>339</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-93.5,259,-93.5,262.5</points>
<connection>
<GID>298</GID>
<name>IN_2</name></connection>
<intersection>262.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-90.5,262.5,-90.5,263</points>
<connection>
<GID>379</GID>
<name>OUT</name></connection>
<intersection>262.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-93.5,262.5,-90.5,262.5</points>
<intersection>-93.5 0</intersection>
<intersection>-90.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>340</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-94.5,259,-94.5,263</points>
<connection>
<GID>298</GID>
<name>IN_3</name></connection>
<connection>
<GID>380</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>358</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-66.5,269,-66.5,274</points>
<connection>
<GID>372</GID>
<name>IN_1</name></connection>
<connection>
<GID>389</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>359</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-70.5,269,-70.5,274</points>
<connection>
<GID>373</GID>
<name>IN_1</name></connection>
<connection>
<GID>388</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>360</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-74.5,269,-74.5,274</points>
<connection>
<GID>374</GID>
<name>IN_1</name></connection>
<connection>
<GID>387</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>361</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-78.5,269,-78.5,274</points>
<connection>
<GID>375</GID>
<name>IN_1</name></connection>
<connection>
<GID>386</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>362</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-83.5,269,-83.5,274</points>
<connection>
<GID>377</GID>
<name>IN_1</name></connection>
<connection>
<GID>385</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>363</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-87.5,269,-87.5,274</points>
<connection>
<GID>378</GID>
<name>IN_1</name></connection>
<connection>
<GID>384</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>364</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-95.5,269,-95.5,274</points>
<connection>
<GID>380</GID>
<name>IN_1</name></connection>
<connection>
<GID>382</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>365</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-91.5,269,-91.5,274</points>
<connection>
<GID>379</GID>
<name>IN_1</name></connection>
<connection>
<GID>383</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>366</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-55,248,-55,282</points>
<intersection>248 1</intersection>
<intersection>282 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-56,248,-50.5,248</points>
<connection>
<GID>307</GID>
<name>OUT_0</name></connection>
<connection>
<GID>319</GID>
<name>N_in0</name></connection>
<intersection>-55 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-67.5,282,-55,282</points>
<intersection>-67.5 3</intersection>
<intersection>-55 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-67.5,280,-67.5,282</points>
<connection>
<GID>389</GID>
<name>IN_1</name></connection>
<intersection>282 2</intersection></vsegment></shape></wire>
<wire>
<ID>367</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-54.5,239,-54.5,282.5</points>
<intersection>239 1</intersection>
<intersection>282.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-56,239,-50.5,239</points>
<connection>
<GID>305</GID>
<name>OUT_0</name></connection>
<connection>
<GID>320</GID>
<name>N_in0</name></connection>
<intersection>-54.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-71.5,282.5,-54.5,282.5</points>
<intersection>-71.5 3</intersection>
<intersection>-54.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-71.5,280,-71.5,282.5</points>
<connection>
<GID>388</GID>
<name>IN_1</name></connection>
<intersection>282.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>368</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-54,230,-54,283</points>
<intersection>230 1</intersection>
<intersection>283 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-56,230,-50.5,230</points>
<connection>
<GID>306</GID>
<name>OUT_0</name></connection>
<connection>
<GID>321</GID>
<name>N_in0</name></connection>
<intersection>-54 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-75.5,283,-54,283</points>
<intersection>-75.5 3</intersection>
<intersection>-54 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-75.5,280,-75.5,283</points>
<connection>
<GID>387</GID>
<name>IN_1</name></connection>
<intersection>283 2</intersection></vsegment></shape></wire>
<wire>
<ID>369</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-53.5,221,-53.5,283.5</points>
<intersection>221 1</intersection>
<intersection>283.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-56,221,-50.5,221</points>
<connection>
<GID>308</GID>
<name>OUT_0</name></connection>
<connection>
<GID>322</GID>
<name>N_in0</name></connection>
<intersection>-53.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-79.5,283.5,-53.5,283.5</points>
<intersection>-79.5 3</intersection>
<intersection>-53.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-79.5,280,-79.5,283.5</points>
<connection>
<GID>386</GID>
<name>IN_1</name></connection>
<intersection>283.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>370</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-53,212,-53,284</points>
<intersection>212 1</intersection>
<intersection>284 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-56,212,-50.5,212</points>
<connection>
<GID>311</GID>
<name>OUT_0</name></connection>
<connection>
<GID>323</GID>
<name>N_in0</name></connection>
<intersection>-53 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-84.5,284,-53,284</points>
<intersection>-84.5 3</intersection>
<intersection>-53 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-84.5,280,-84.5,284</points>
<connection>
<GID>385</GID>
<name>IN_1</name></connection>
<intersection>284 2</intersection></vsegment></shape></wire>
<wire>
<ID>371</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-52.5,203,-52.5,284.5</points>
<intersection>203 1</intersection>
<intersection>284.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-56,203,-50.5,203</points>
<connection>
<GID>324</GID>
<name>N_in0</name></connection>
<connection>
<GID>309</GID>
<name>OUT_0</name></connection>
<intersection>-52.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-88.5,284.5,-52.5,284.5</points>
<intersection>-88.5 3</intersection>
<intersection>-52.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-88.5,280,-88.5,284.5</points>
<connection>
<GID>384</GID>
<name>IN_1</name></connection>
<intersection>284.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>372</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-52,194,-52,285</points>
<intersection>194 1</intersection>
<intersection>285 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-56,194,-50.5,194</points>
<connection>
<GID>310</GID>
<name>OUT_0</name></connection>
<connection>
<GID>325</GID>
<name>N_in0</name></connection>
<intersection>-52 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-92.5,285,-52,285</points>
<intersection>-92.5 3</intersection>
<intersection>-52 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-92.5,280,-92.5,285</points>
<connection>
<GID>383</GID>
<name>IN_1</name></connection>
<intersection>285 2</intersection></vsegment></shape></wire>
<wire>
<ID>373</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-51.5,185,-51.5,285.5</points>
<intersection>185 1</intersection>
<intersection>285.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-56,185,-50.5,185</points>
<connection>
<GID>312</GID>
<name>OUT_0</name></connection>
<connection>
<GID>326</GID>
<name>N_in0</name></connection>
<intersection>-51.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-96.5,285.5,-51.5,285.5</points>
<intersection>-96.5 3</intersection>
<intersection>-51.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-96.5,280,-96.5,285.5</points>
<connection>
<GID>382</GID>
<name>IN_1</name></connection>
<intersection>285.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>375</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-94.5,280,-94.5,281</points>
<connection>
<GID>382</GID>
<name>IN_0</name></connection>
<intersection>281 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-26,249.5,-26,281</points>
<intersection>249.5 10</intersection>
<intersection>281 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-94.5,281,-26,281</points>
<intersection>-94.5 0</intersection>
<intersection>-90.5 3</intersection>
<intersection>-86.5 4</intersection>
<intersection>-82.5 5</intersection>
<intersection>-77.5 6</intersection>
<intersection>-73.5 7</intersection>
<intersection>-69.5 8</intersection>
<intersection>-65.5 9</intersection>
<intersection>-26 1</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-90.5,280,-90.5,281</points>
<connection>
<GID>383</GID>
<name>IN_0</name></connection>
<intersection>281 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-86.5,280,-86.5,281</points>
<connection>
<GID>384</GID>
<name>IN_0</name></connection>
<intersection>281 2</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-82.5,280,-82.5,281</points>
<connection>
<GID>385</GID>
<name>IN_0</name></connection>
<intersection>281 2</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-77.5,280,-77.5,281</points>
<connection>
<GID>386</GID>
<name>IN_0</name></connection>
<intersection>281 2</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>-73.5,280,-73.5,281</points>
<connection>
<GID>387</GID>
<name>IN_0</name></connection>
<intersection>281 2</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>-69.5,280,-69.5,281</points>
<connection>
<GID>388</GID>
<name>IN_0</name></connection>
<intersection>281 2</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>-65.5,280,-65.5,281</points>
<connection>
<GID>389</GID>
<name>IN_0</name></connection>
<intersection>281 2</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-26,249.5,37,249.5</points>
<intersection>-26 1</intersection>
<intersection>37 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>37,232.5,37,249.5</points>
<connection>
<GID>393</GID>
<name>OUT_0</name></connection>
<intersection>249.5 10</intersection></vsegment></shape></wire>
<wire>
<ID>387</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,306.5,32,312.5</points>
<intersection>306.5 3</intersection>
<intersection>312.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>30,312.5,32,312.5</points>
<connection>
<GID>408</GID>
<name>OUT</name></connection>
<intersection>30 8</intersection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>32,306.5,33,306.5</points>
<connection>
<GID>409</GID>
<name>IN_0</name></connection>
<intersection>32 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>30,312.5,30,313</points>
<connection>
<GID>417</GID>
<name>N_in0</name></connection>
<intersection>312.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>388</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,306.5,32,312.5</points>
<intersection>306.5 5</intersection>
<intersection>312.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>32,312.5,34,312.5</points>
<connection>
<GID>409</GID>
<name>OUT</name></connection>
<intersection>32 0</intersection>
<intersection>34 10</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>31,306.5,32,306.5</points>
<connection>
<GID>408</GID>
<name>IN_1</name></connection>
<intersection>32 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>34,312.5,34,313</points>
<connection>
<GID>419</GID>
<name>N_in0</name></connection>
<intersection>312.5 2</intersection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>-1.20056,382.685,1136.8,-478.315</PageViewport>
<gate>
<ID>89</ID>
<type>AF_DFF_LOW</type>
<position>47,-21.5</position>
<input>
<ID>IN_0</ID>111 </input>
<output>
<ID>OUT_0</ID>107 </output>
<input>
<ID>clear</ID>101 </input>
<input>
<ID>clock</ID>116 </input>
<input>
<ID>clock_enable</ID>117 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>90</ID>
<type>AF_DFF_LOW</type>
<position>47,-30</position>
<input>
<ID>IN_0</ID>112 </input>
<output>
<ID>OUT_0</ID>108 </output>
<input>
<ID>clear</ID>102 </input>
<input>
<ID>clock</ID>116 </input>
<input>
<ID>clock_enable</ID>117 </input>
<input>
<ID>set</ID>101 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>91</ID>
<type>AF_DFF_LOW</type>
<position>47,-38.5</position>
<input>
<ID>IN_0</ID>113 </input>
<output>
<ID>OUT_0</ID>109 </output>
<input>
<ID>clear</ID>103 </input>
<input>
<ID>clock</ID>116 </input>
<input>
<ID>clock_enable</ID>117 </input>
<input>
<ID>set</ID>102 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>92</ID>
<type>AF_DFF_LOW</type>
<position>47,-47</position>
<input>
<ID>IN_0</ID>114 </input>
<output>
<ID>OUT_0</ID>110 </output>
<input>
<ID>clear</ID>122 </input>
<input>
<ID>clock</ID>116 </input>
<input>
<ID>clock_enable</ID>117 </input>
<input>
<ID>set</ID>103 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>93</ID>
<type>AF_DFF_LOW</type>
<position>60.5,-21.5</position>
<input>
<ID>IN_0</ID>107 </input>
<output>
<ID>OUT_0</ID>135 </output>
<input>
<ID>clear</ID>104 </input>
<input>
<ID>clock</ID>117 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>94</ID>
<type>AF_DFF_LOW</type>
<position>60.5,-30</position>
<input>
<ID>IN_0</ID>108 </input>
<output>
<ID>OUT_0</ID>136 </output>
<input>
<ID>clear</ID>105 </input>
<input>
<ID>clock</ID>117 </input>
<input>
<ID>set</ID>104 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>95</ID>
<type>AF_DFF_LOW</type>
<position>60.5,-38.5</position>
<input>
<ID>IN_0</ID>109 </input>
<output>
<ID>OUT_0</ID>137 </output>
<input>
<ID>clear</ID>106 </input>
<input>
<ID>clock</ID>117 </input>
<input>
<ID>set</ID>105 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>96</ID>
<type>AF_DFF_LOW</type>
<position>60.5,-47</position>
<input>
<ID>IN_0</ID>110 </input>
<output>
<ID>OUT_0</ID>138 </output>
<input>
<ID>clear</ID>130 </input>
<input>
<ID>clock</ID>117 </input>
<input>
<ID>set</ID>106 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>97</ID>
<type>AE_FULLADDER_4BIT</type>
<position>31,-43.5</position>
<input>
<ID>IN_0</ID>135 </input>
<input>
<ID>IN_1</ID>136 </input>
<input>
<ID>IN_2</ID>137 </input>
<input>
<ID>IN_3</ID>138 </input>
<input>
<ID>IN_B_0</ID>115 </input>
<output>
<ID>OUT_0</ID>111 </output>
<output>
<ID>OUT_1</ID>112 </output>
<output>
<ID>OUT_2</ID>113 </output>
<output>
<ID>OUT_3</ID>114 </output>
<output>
<ID>carry_out</ID>118 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>98</ID>
<type>DA_FROM</type>
<position>37,-7</position>
<input>
<ID>IN_0</ID>116 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>99</ID>
<type>AA_TOGGLE</type>
<position>24,-38.5</position>
<output>
<ID>OUT_0</ID>115 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>100</ID>
<type>DA_FROM</type>
<position>37,-9</position>
<input>
<ID>IN_0</ID>117 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID nclk</lparam></gate>
<gate>
<ID>101</ID>
<type>AE_FULLADDER_4BIT</type>
<position>31,-60.5</position>
<input>
<ID>IN_0</ID>139 </input>
<input>
<ID>IN_1</ID>140 </input>
<input>
<ID>IN_2</ID>141 </input>
<input>
<ID>IN_3</ID>142 </input>
<output>
<ID>OUT_0</ID>123 </output>
<output>
<ID>OUT_1</ID>124 </output>
<output>
<ID>OUT_2</ID>125 </output>
<output>
<ID>OUT_3</ID>126 </output>
<input>
<ID>carry_in</ID>118 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>102</ID>
<type>AF_DFF_LOW</type>
<position>47,-57</position>
<input>
<ID>IN_0</ID>123 </input>
<output>
<ID>OUT_0</ID>131 </output>
<input>
<ID>clear</ID>119 </input>
<input>
<ID>clock</ID>116 </input>
<input>
<ID>clock_enable</ID>117 </input>
<input>
<ID>set</ID>122 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>103</ID>
<type>AF_DFF_LOW</type>
<position>47,-65.5</position>
<input>
<ID>IN_0</ID>124 </input>
<output>
<ID>OUT_0</ID>132 </output>
<input>
<ID>clear</ID>120 </input>
<input>
<ID>clock</ID>116 </input>
<input>
<ID>clock_enable</ID>117 </input>
<input>
<ID>set</ID>119 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>104</ID>
<type>AF_DFF_LOW</type>
<position>47,-74</position>
<input>
<ID>IN_0</ID>125 </input>
<output>
<ID>OUT_0</ID>133 </output>
<input>
<ID>clear</ID>121 </input>
<input>
<ID>clock</ID>116 </input>
<input>
<ID>clock_enable</ID>117 </input>
<input>
<ID>set</ID>120 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>105</ID>
<type>AF_DFF_LOW</type>
<position>47,-82.5</position>
<input>
<ID>IN_0</ID>126 </input>
<output>
<ID>OUT_0</ID>134 </output>
<input>
<ID>clock</ID>116 </input>
<input>
<ID>clock_enable</ID>117 </input>
<input>
<ID>set</ID>121 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>106</ID>
<type>AF_DFF_LOW</type>
<position>60.5,-57</position>
<input>
<ID>IN_0</ID>131 </input>
<output>
<ID>OUT_0</ID>139 </output>
<input>
<ID>clear</ID>127 </input>
<input>
<ID>clock</ID>117 </input>
<input>
<ID>set</ID>130 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>107</ID>
<type>AF_DFF_LOW</type>
<position>60.5,-65.5</position>
<input>
<ID>IN_0</ID>132 </input>
<output>
<ID>OUT_0</ID>140 </output>
<input>
<ID>clear</ID>128 </input>
<input>
<ID>clock</ID>117 </input>
<input>
<ID>set</ID>127 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>108</ID>
<type>AF_DFF_LOW</type>
<position>60.5,-74</position>
<input>
<ID>IN_0</ID>133 </input>
<output>
<ID>OUT_0</ID>141 </output>
<input>
<ID>clear</ID>129 </input>
<input>
<ID>clock</ID>117 </input>
<input>
<ID>set</ID>128 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>109</ID>
<type>AF_DFF_LOW</type>
<position>60.5,-82.5</position>
<input>
<ID>IN_0</ID>134 </input>
<output>
<ID>OUT_0</ID>142 </output>
<input>
<ID>clock</ID>117 </input>
<input>
<ID>set</ID>129 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>110</ID>
<type>HA_JUNC_2</type>
<position>73,-19.5</position>
<input>
<ID>N_in0</ID>135 </input>
<input>
<ID>N_in1</ID>150 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>111</ID>
<type>HA_JUNC_2</type>
<position>73,-28</position>
<input>
<ID>N_in0</ID>136 </input>
<input>
<ID>N_in1</ID>149 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>112</ID>
<type>HA_JUNC_2</type>
<position>73,-36.5</position>
<input>
<ID>N_in0</ID>137 </input>
<input>
<ID>N_in1</ID>148 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>113</ID>
<type>HA_JUNC_2</type>
<position>73,-45</position>
<input>
<ID>N_in0</ID>138 </input>
<input>
<ID>N_in1</ID>147 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>114</ID>
<type>HA_JUNC_2</type>
<position>73,-55</position>
<input>
<ID>N_in0</ID>139 </input>
<input>
<ID>N_in1</ID>146 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>115</ID>
<type>HA_JUNC_2</type>
<position>73,-63.5</position>
<input>
<ID>N_in0</ID>140 </input>
<input>
<ID>N_in1</ID>145 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>116</ID>
<type>HA_JUNC_2</type>
<position>73,-72</position>
<input>
<ID>N_in0</ID>141 </input>
<input>
<ID>N_in1</ID>144 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>117</ID>
<type>HA_JUNC_2</type>
<position>73.5,-80.5</position>
<input>
<ID>N_in0</ID>142 </input>
<input>
<ID>N_in1</ID>143 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>118</ID>
<type>BE_ROM_8x8</type>
<position>100,-84</position>
<input>
<ID>ADDRESS_0</ID>150 </input>
<input>
<ID>ADDRESS_1</ID>149 </input>
<input>
<ID>ADDRESS_2</ID>148 </input>
<input>
<ID>ADDRESS_3</ID>147 </input>
<input>
<ID>ADDRESS_4</ID>146 </input>
<input>
<ID>ADDRESS_5</ID>145 </input>
<input>
<ID>ADDRESS_6</ID>144 </input>
<input>
<ID>ADDRESS_7</ID>143 </input>
<input>
<ID>ENABLE_0</ID>151 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam></gate>
<gate>
<ID>119</ID>
<type>AA_TOGGLE</type>
<position>108,-84.5</position>
<output>
<ID>OUT_0</ID>151 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>120</ID>
<type>AO_XNOR2</type>
<position>23,42.5</position>
<input>
<ID>IN_0</ID>152 </input>
<input>
<ID>IN_1</ID>159 </input>
<output>
<ID>OUT</ID>169 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>121</ID>
<type>AO_XNOR2</type>
<position>27,42.5</position>
<input>
<ID>IN_0</ID>153 </input>
<input>
<ID>IN_1</ID>160 </input>
<output>
<ID>OUT</ID>167 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>122</ID>
<type>AO_XNOR2</type>
<position>31,42.5</position>
<input>
<ID>IN_0</ID>154 </input>
<input>
<ID>IN_1</ID>161 </input>
<output>
<ID>OUT</ID>168 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>123</ID>
<type>AO_XNOR2</type>
<position>35,42.5</position>
<input>
<ID>IN_0</ID>155 </input>
<input>
<ID>IN_1</ID>162 </input>
<output>
<ID>OUT</ID>170 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>124</ID>
<type>HA_JUNC_2</type>
<position>20,38.5</position>
<input>
<ID>N_in1</ID>152 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>125</ID>
<type>HA_JUNC_2</type>
<position>20,37.5</position>
<input>
<ID>N_in1</ID>153 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>126</ID>
<type>HA_JUNC_2</type>
<position>20,36.5</position>
<input>
<ID>N_in1</ID>154 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>127</ID>
<type>HA_JUNC_2</type>
<position>20,35.5</position>
<input>
<ID>N_in1</ID>155 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>128</ID>
<type>HA_JUNC_2</type>
<position>20,34.5</position>
<input>
<ID>N_in1</ID>156 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>129</ID>
<type>HA_JUNC_2</type>
<position>20,33.5</position>
<input>
<ID>N_in1</ID>183 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>130</ID>
<type>HA_JUNC_2</type>
<position>20,32.5</position>
<input>
<ID>N_in1</ID>157 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>131</ID>
<type>HA_JUNC_2</type>
<position>20,31.5</position>
<input>
<ID>N_in1</ID>158 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>132</ID>
<type>AO_XNOR2</type>
<position>39,42.5</position>
<input>
<ID>IN_0</ID>156 </input>
<input>
<ID>IN_1</ID>163 </input>
<output>
<ID>OUT</ID>173 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>133</ID>
<type>AO_XNOR2</type>
<position>43,42.5</position>
<input>
<ID>IN_0</ID>183 </input>
<input>
<ID>IN_1</ID>164 </input>
<output>
<ID>OUT</ID>171 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>134</ID>
<type>AO_XNOR2</type>
<position>47,42.5</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>165 </input>
<output>
<ID>OUT</ID>172 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>135</ID>
<type>AO_XNOR2</type>
<position>51,42.5</position>
<input>
<ID>IN_0</ID>158 </input>
<input>
<ID>IN_1</ID>166 </input>
<output>
<ID>OUT</ID>185 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>136</ID>
<type>HA_JUNC_2</type>
<position>20,26.5</position>
<input>
<ID>N_in1</ID>159 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>137</ID>
<type>HA_JUNC_2</type>
<position>20,25.5</position>
<input>
<ID>N_in1</ID>160 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>138</ID>
<type>HA_JUNC_2</type>
<position>20,24.5</position>
<input>
<ID>N_in1</ID>161 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>139</ID>
<type>HA_JUNC_2</type>
<position>20,23.5</position>
<input>
<ID>N_in1</ID>162 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>140</ID>
<type>HA_JUNC_2</type>
<position>20,22.5</position>
<input>
<ID>N_in1</ID>163 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>141</ID>
<type>HA_JUNC_2</type>
<position>20,21.5</position>
<input>
<ID>N_in1</ID>164 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>142</ID>
<type>HA_JUNC_2</type>
<position>20,20.5</position>
<input>
<ID>N_in1</ID>165 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>143</ID>
<type>HA_JUNC_2</type>
<position>20,19.5</position>
<input>
<ID>N_in1</ID>166 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>144</ID>
<type>AA_AND4</type>
<position>10,57.5</position>
<input>
<ID>IN_0</ID>169 </input>
<input>
<ID>IN_1</ID>167 </input>
<input>
<ID>IN_2</ID>168 </input>
<input>
<ID>IN_3</ID>170 </input>
<output>
<ID>OUT</ID>174 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>145</ID>
<type>AA_AND4</type>
<position>18,57.5</position>
<input>
<ID>IN_0</ID>173 </input>
<input>
<ID>IN_1</ID>171 </input>
<input>
<ID>IN_2</ID>172 </input>
<input>
<ID>IN_3</ID>185 </input>
<output>
<ID>OUT</ID>175 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>146</ID>
<type>AA_AND2</type>
<position>14,65.5</position>
<input>
<ID>IN_0</ID>174 </input>
<input>
<ID>IN_1</ID>175 </input>
<output>
<ID>OUT</ID>198 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>147</ID>
<type>AA_AND2</type>
<position>56,58.5</position>
<input>
<ID>IN_0</ID>152 </input>
<input>
<ID>IN_1</ID>176 </input>
<output>
<ID>OUT</ID>190 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>148</ID>
<type>AE_SMALL_INVERTER</type>
<position>57,41.5</position>
<input>
<ID>IN_0</ID>159 </input>
<output>
<ID>OUT_0</ID>176 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>149</ID>
<type>AA_AND3</type>
<position>62,58.5</position>
<input>
<ID>IN_0</ID>169 </input>
<input>
<ID>IN_1</ID>153 </input>
<input>
<ID>IN_2</ID>177 </input>
<output>
<ID>OUT</ID>191 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>150</ID>
<type>AE_SMALL_INVERTER</type>
<position>64,41.5</position>
<input>
<ID>IN_0</ID>160 </input>
<output>
<ID>OUT_0</ID>177 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>151</ID>
<type>AA_AND4</type>
<position>70,58.5</position>
<input>
<ID>IN_0</ID>169 </input>
<input>
<ID>IN_1</ID>167 </input>
<input>
<ID>IN_2</ID>154 </input>
<input>
<ID>IN_3</ID>178 </input>
<output>
<ID>OUT</ID>192 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>152</ID>
<type>AE_SMALL_INVERTER</type>
<position>73,41.5</position>
<input>
<ID>IN_0</ID>161 </input>
<output>
<ID>OUT_0</ID>178 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>153</ID>
<type>AA_AND3</type>
<position>78,58.5</position>
<input>
<ID>IN_0</ID>169 </input>
<input>
<ID>IN_1</ID>167 </input>
<input>
<ID>IN_2</ID>168 </input>
<output>
<ID>OUT</ID>179 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>154</ID>
<type>AA_AND3</type>
<position>86,58.5</position>
<input>
<ID>IN_0</ID>179 </input>
<input>
<ID>IN_1</ID>155 </input>
<input>
<ID>IN_2</ID>180 </input>
<output>
<ID>OUT</ID>193 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>155</ID>
<type>AE_SMALL_INVERTER</type>
<position>88,41.5</position>
<input>
<ID>IN_0</ID>162 </input>
<output>
<ID>OUT_0</ID>180 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>156</ID>
<type>AA_AND4</type>
<position>94,58.5</position>
<input>
<ID>IN_0</ID>169 </input>
<input>
<ID>IN_1</ID>167 </input>
<input>
<ID>IN_2</ID>168 </input>
<input>
<ID>IN_3</ID>170 </input>
<output>
<ID>OUT</ID>181 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>157</ID>
<type>AA_AND3</type>
<position>103,58.5</position>
<input>
<ID>IN_0</ID>181 </input>
<input>
<ID>IN_1</ID>156 </input>
<input>
<ID>IN_2</ID>182 </input>
<output>
<ID>OUT</ID>194 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>158</ID>
<type>AE_SMALL_INVERTER</type>
<position>105,41.5</position>
<input>
<ID>IN_0</ID>163 </input>
<output>
<ID>OUT_0</ID>182 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>159</ID>
<type>AA_AND4</type>
<position>111,58.5</position>
<input>
<ID>IN_0</ID>169 </input>
<input>
<ID>IN_1</ID>167 </input>
<input>
<ID>IN_2</ID>168 </input>
<input>
<ID>IN_3</ID>170 </input>
<output>
<ID>OUT</ID>184 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>160</ID>
<type>AA_AND4</type>
<position>121,58.5</position>
<input>
<ID>IN_0</ID>184 </input>
<input>
<ID>IN_1</ID>173 </input>
<input>
<ID>IN_2</ID>183 </input>
<input>
<ID>IN_3</ID>188 </input>
<output>
<ID>OUT</ID>195 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>161</ID>
<type>DA_AND8</type>
<position>139,58.5</position>
<input>
<ID>IN_0</ID>169 </input>
<input>
<ID>IN_1</ID>167 </input>
<input>
<ID>IN_2</ID>168 </input>
<input>
<ID>IN_3</ID>170 </input>
<input>
<ID>IN_4</ID>173 </input>
<input>
<ID>IN_5</ID>171 </input>
<input>
<ID>IN_6</ID>172 </input>
<input>
<ID>IN_7</ID>158 </input>
<output>
<ID>OUT</ID>186 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>162</ID>
<type>AA_AND2</type>
<position>147,58.5</position>
<input>
<ID>IN_0</ID>186 </input>
<input>
<ID>IN_1</ID>187 </input>
<output>
<ID>OUT</ID>197 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>163</ID>
<type>AE_SMALL_INVERTER</type>
<position>148,41.5</position>
<input>
<ID>IN_0</ID>166 </input>
<output>
<ID>OUT_0</ID>187 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>164</ID>
<type>AE_SMALL_INVERTER</type>
<position>124,41.5</position>
<input>
<ID>IN_0</ID>164 </input>
<output>
<ID>OUT_0</ID>188 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>165</ID>
<type>DA_AND8</type>
<position>130,58.5</position>
<input>
<ID>IN_0</ID>169 </input>
<input>
<ID>IN_1</ID>167 </input>
<input>
<ID>IN_2</ID>168 </input>
<input>
<ID>IN_3</ID>170 </input>
<input>
<ID>IN_4</ID>173 </input>
<input>
<ID>IN_5</ID>171 </input>
<input>
<ID>IN_6</ID>157 </input>
<input>
<ID>IN_7</ID>189 </input>
<output>
<ID>OUT</ID>196 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>166</ID>
<type>AE_SMALL_INVERTER</type>
<position>133.5,41.5</position>
<input>
<ID>IN_0</ID>165 </input>
<output>
<ID>OUT_0</ID>189 </output>
<gparam>angle 90</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>167</ID>
<type>DE_OR8</type>
<position>50,73.5</position>
<input>
<ID>IN_0</ID>190 </input>
<input>
<ID>IN_1</ID>191 </input>
<input>
<ID>IN_2</ID>192 </input>
<input>
<ID>IN_3</ID>193 </input>
<input>
<ID>IN_4</ID>197 </input>
<input>
<ID>IN_5</ID>196 </input>
<input>
<ID>IN_6</ID>195 </input>
<input>
<ID>IN_7</ID>194 </input>
<output>
<ID>OUT</ID>199 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>168</ID>
<type>BE_NOR2</type>
<position>30.5,73.5</position>
<input>
<ID>IN_0</ID>198 </input>
<input>
<ID>IN_1</ID>199 </input>
<output>
<ID>OUT</ID>200 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>169</ID>
<type>HA_JUNC_2</type>
<position>50,80.5</position>
<input>
<ID>N_in0</ID>199 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>170</ID>
<type>HA_JUNC_2</type>
<position>30.5,80.5</position>
<input>
<ID>N_in0</ID>200 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>171</ID>
<type>HA_JUNC_2</type>
<position>14,80.5</position>
<input>
<ID>N_in0</ID>198 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 90</gparam></gate>
<gate>
<ID>172</ID>
<type>AA_LABEL</type>
<position>17.5,35.5</position>
<gparam>LABEL_TEXT a</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>173</ID>
<type>AA_LABEL</type>
<position>17.5,24</position>
<gparam>LABEL_TEXT b</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>174</ID>
<type>AA_LABEL</type>
<position>18.5,81</position>
<gparam>LABEL_TEXT a = b</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>175</ID>
<type>AA_LABEL</type>
<position>35,81</position>
<gparam>LABEL_TEXT a  b</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>176</ID>
<type>AA_LABEL</type>
<position>54.5,81</position>
<gparam>LABEL_TEXT a > b</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>193</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,65.5,49.5,70.5</points>
<connection>
<GID>167</GID>
<name>IN_3</name></connection>
<intersection>65.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>86,61.5,86,65.5</points>
<connection>
<GID>154</GID>
<name>OUT</name></connection>
<intersection>65.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>49.5,65.5,86,65.5</points>
<intersection>49.5 0</intersection>
<intersection>86 1</intersection></hsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,66.5,50.5,70.5</points>
<connection>
<GID>167</GID>
<name>IN_7</name></connection>
<intersection>66.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>103,61.5,103,66.5</points>
<connection>
<GID>157</GID>
<name>OUT</name></connection>
<intersection>66.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>50.5,66.5,103,66.5</points>
<intersection>50.5 0</intersection>
<intersection>103 1</intersection></hsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,67.5,51.5,70.5</points>
<connection>
<GID>167</GID>
<name>IN_6</name></connection>
<intersection>67.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>121,61.5,121,67.5</points>
<connection>
<GID>160</GID>
<name>OUT</name></connection>
<intersection>67.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>51.5,67.5,121,67.5</points>
<intersection>51.5 0</intersection>
<intersection>121 1</intersection></hsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,68.5,52.5,70.5</points>
<connection>
<GID>167</GID>
<name>IN_5</name></connection>
<intersection>68.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>130,61.5,130,68.5</points>
<connection>
<GID>165</GID>
<name>OUT</name></connection>
<intersection>68.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>52.5,68.5,130,68.5</points>
<intersection>52.5 0</intersection>
<intersection>130 1</intersection></hsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,69.5,53.5,70.5</points>
<connection>
<GID>167</GID>
<name>IN_4</name></connection>
<intersection>69.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>147,61.5,147,69.5</points>
<connection>
<GID>162</GID>
<name>OUT</name></connection>
<intersection>69.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>53.5,69.5,147,69.5</points>
<intersection>53.5 0</intersection>
<intersection>147 1</intersection></hsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14,68.5,14,79.5</points>
<connection>
<GID>171</GID>
<name>N_in0</name></connection>
<connection>
<GID>146</GID>
<name>OUT</name></connection>
<intersection>69.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>29.5,69.5,29.5,70.5</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<intersection>69.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>14,69.5,29.5,69.5</points>
<intersection>14 0</intersection>
<intersection>29.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,69.5,31.5,70.5</points>
<connection>
<GID>168</GID>
<name>IN_1</name></connection>
<intersection>69.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>40,69.5,40,78.5</points>
<intersection>69.5 2</intersection>
<intersection>78.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>31.5,69.5,40,69.5</points>
<intersection>31.5 0</intersection>
<intersection>40 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>40,78.5,50,78.5</points>
<intersection>40 1</intersection>
<intersection>50 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>50,77.5,50,79.5</points>
<connection>
<GID>169</GID>
<name>N_in0</name></connection>
<connection>
<GID>167</GID>
<name>OUT</name></connection>
<intersection>78.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>30.5,76.5,30.5,79.5</points>
<connection>
<GID>170</GID>
<name>N_in0</name></connection>
<connection>
<GID>168</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-26,47,-25.5</points>
<connection>
<GID>90</GID>
<name>set</name></connection>
<connection>
<GID>89</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-34.5,47,-34</points>
<connection>
<GID>91</GID>
<name>set</name></connection>
<connection>
<GID>90</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-43,47,-42.5</points>
<connection>
<GID>92</GID>
<name>set</name></connection>
<connection>
<GID>91</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-26,60.5,-25.5</points>
<connection>
<GID>94</GID>
<name>set</name></connection>
<connection>
<GID>93</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-34.5,60.5,-34</points>
<connection>
<GID>95</GID>
<name>set</name></connection>
<connection>
<GID>94</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-43,60.5,-42.5</points>
<connection>
<GID>96</GID>
<name>set</name></connection>
<connection>
<GID>95</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-19.5,57.5,-19.5</points>
<connection>
<GID>89</GID>
<name>OUT_0</name></connection>
<connection>
<GID>93</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-28,57.5,-28</points>
<connection>
<GID>90</GID>
<name>OUT_0</name></connection>
<connection>
<GID>94</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-36.5,57.5,-36.5</points>
<connection>
<GID>91</GID>
<name>OUT_0</name></connection>
<connection>
<GID>95</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-45,57.5,-45</points>
<connection>
<GID>92</GID>
<name>OUT_0</name></connection>
<connection>
<GID>96</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-42,36,-19.5</points>
<intersection>-42 2</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-19.5,44,-19.5</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35,-42,36,-42</points>
<connection>
<GID>97</GID>
<name>OUT_0</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-43,37,-28</points>
<intersection>-43 2</intersection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,-28,44,-28</points>
<connection>
<GID>90</GID>
<name>IN_0</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35,-43,37,-43</points>
<connection>
<GID>97</GID>
<name>OUT_1</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35,-44,38,-44</points>
<connection>
<GID>97</GID>
<name>OUT_2</name></connection>
<intersection>38 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>38,-44,38,-36.5</points>
<intersection>-44 1</intersection>
<intersection>-36.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>38,-36.5,44,-36.5</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<intersection>38 4</intersection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35,-45,44,-45</points>
<connection>
<GID>97</GID>
<name>OUT_3</name></connection>
<connection>
<GID>92</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>26,-38.5,27,-38.5</points>
<connection>
<GID>99</GID>
<name>OUT_0</name></connection>
<connection>
<GID>97</GID>
<name>IN_B_0</name></connection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,-82.5,41,-7</points>
<intersection>-82.5 10</intersection>
<intersection>-74 13</intersection>
<intersection>-65.5 12</intersection>
<intersection>-57 11</intersection>
<intersection>-47 8</intersection>
<intersection>-38.5 6</intersection>
<intersection>-30 4</intersection>
<intersection>-21.5 1</intersection>
<intersection>-7 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41,-21.5,44,-21.5</points>
<connection>
<GID>89</GID>
<name>clock</name></connection>
<intersection>41 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>39,-7,41,-7</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>41 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>41,-30,44,-30</points>
<connection>
<GID>90</GID>
<name>clock</name></connection>
<intersection>41 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>41,-38.5,44,-38.5</points>
<connection>
<GID>91</GID>
<name>clock</name></connection>
<intersection>41 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>41,-47,44,-47</points>
<connection>
<GID>92</GID>
<name>clock</name></connection>
<intersection>41 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>41,-82.5,44,-82.5</points>
<connection>
<GID>105</GID>
<name>clock</name></connection>
<intersection>41 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>41,-57,44,-57</points>
<connection>
<GID>102</GID>
<name>clock</name></connection>
<intersection>41 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>41,-65.5,44,-65.5</points>
<connection>
<GID>103</GID>
<name>clock</name></connection>
<intersection>41 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>41,-74,44,-74</points>
<connection>
<GID>104</GID>
<name>clock</name></connection>
<intersection>41 0</intersection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-84.5,40,-9</points>
<intersection>-84.5 23</intersection>
<intersection>-76 16</intersection>
<intersection>-67.5 17</intersection>
<intersection>-59 18</intersection>
<intersection>-49 9</intersection>
<intersection>-40.5 5</intersection>
<intersection>-32 6</intersection>
<intersection>-23.5 1</intersection>
<intersection>-9 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-23.5,44,-23.5</points>
<connection>
<GID>89</GID>
<name>clock_enable</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>39,-9,55.5,-9</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>40 0</intersection>
<intersection>55.5 7</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>40,-40.5,44,-40.5</points>
<connection>
<GID>91</GID>
<name>clock_enable</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>40,-32,44,-32</points>
<connection>
<GID>90</GID>
<name>clock_enable</name></connection>
<intersection>40 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>55.5,-82.5,55.5,-9</points>
<intersection>-82.5 24</intersection>
<intersection>-74 27</intersection>
<intersection>-65.5 26</intersection>
<intersection>-57 25</intersection>
<intersection>-47 10</intersection>
<intersection>-38.5 11</intersection>
<intersection>-30 12</intersection>
<intersection>-21.5 13</intersection>
<intersection>-9 2</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>40,-49,44,-49</points>
<connection>
<GID>92</GID>
<name>clock_enable</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>55.5,-47,57.5,-47</points>
<connection>
<GID>96</GID>
<name>clock</name></connection>
<intersection>55.5 7</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>55.5,-38.5,57.5,-38.5</points>
<connection>
<GID>95</GID>
<name>clock</name></connection>
<intersection>55.5 7</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>55.5,-30,57.5,-30</points>
<connection>
<GID>94</GID>
<name>clock</name></connection>
<intersection>55.5 7</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>55.5,-21.5,57.5,-21.5</points>
<connection>
<GID>93</GID>
<name>clock</name></connection>
<intersection>55.5 7</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>40,-76,44,-76</points>
<connection>
<GID>104</GID>
<name>clock_enable</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>40,-67.5,44,-67.5</points>
<connection>
<GID>103</GID>
<name>clock_enable</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>40,-59,44,-59</points>
<connection>
<GID>102</GID>
<name>clock_enable</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>40,-84.5,44,-84.5</points>
<connection>
<GID>105</GID>
<name>clock_enable</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>55.5,-82.5,57.5,-82.5</points>
<connection>
<GID>109</GID>
<name>clock</name></connection>
<intersection>55.5 7</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>55.5,-57,57.5,-57</points>
<connection>
<GID>106</GID>
<name>clock</name></connection>
<intersection>55.5 7</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>55.5,-65.5,57.5,-65.5</points>
<connection>
<GID>107</GID>
<name>clock</name></connection>
<intersection>55.5 7</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>55.5,-74,57.5,-74</points>
<connection>
<GID>108</GID>
<name>clock</name></connection>
<intersection>55.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-52.5,30,-51.5</points>
<connection>
<GID>101</GID>
<name>carry_in</name></connection>
<connection>
<GID>97</GID>
<name>carry_out</name></connection></vsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-61.5,47,-61</points>
<connection>
<GID>103</GID>
<name>set</name></connection>
<connection>
<GID>102</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-70,47,-69.5</points>
<connection>
<GID>104</GID>
<name>set</name></connection>
<connection>
<GID>103</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-78.5,47,-78</points>
<connection>
<GID>105</GID>
<name>set</name></connection>
<connection>
<GID>104</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-53,47,-51</points>
<connection>
<GID>102</GID>
<name>set</name></connection>
<connection>
<GID>92</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-59,36,-55</points>
<intersection>-59 2</intersection>
<intersection>-55 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-55,44,-55</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35,-59,36,-59</points>
<connection>
<GID>101</GID>
<name>OUT_0</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-63.5,38,-60</points>
<intersection>-63.5 1</intersection>
<intersection>-60 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38,-63.5,44,-63.5</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35,-60,38,-60</points>
<connection>
<GID>101</GID>
<name>OUT_1</name></connection>
<intersection>38 0</intersection></hsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-72,37,-61</points>
<intersection>-72 1</intersection>
<intersection>-61 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,-72,44,-72</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35,-61,37,-61</points>
<connection>
<GID>101</GID>
<name>OUT_2</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-80.5,36,-62</points>
<intersection>-80.5 1</intersection>
<intersection>-62 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-80.5,44,-80.5</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35,-62,36,-62</points>
<connection>
<GID>101</GID>
<name>OUT_3</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-61.5,60.5,-61</points>
<connection>
<GID>107</GID>
<name>set</name></connection>
<connection>
<GID>106</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-70,60.5,-69.5</points>
<connection>
<GID>108</GID>
<name>set</name></connection>
<connection>
<GID>107</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-78.5,60.5,-78</points>
<connection>
<GID>109</GID>
<name>set</name></connection>
<connection>
<GID>108</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-53,60.5,-51</points>
<connection>
<GID>106</GID>
<name>set</name></connection>
<connection>
<GID>96</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-55,57.5,-55</points>
<connection>
<GID>102</GID>
<name>OUT_0</name></connection>
<connection>
<GID>106</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-63.5,57.5,-63.5</points>
<connection>
<GID>103</GID>
<name>OUT_0</name></connection>
<connection>
<GID>107</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-72,57.5,-72</points>
<connection>
<GID>104</GID>
<name>OUT_0</name></connection>
<connection>
<GID>108</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50,-80.5,57.5,-80.5</points>
<connection>
<GID>105</GID>
<name>OUT_0</name></connection>
<connection>
<GID>109</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,-94,19,-45.5</points>
<intersection>-94 2</intersection>
<intersection>-45.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19,-45.5,27,-45.5</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>19 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>19,-94,71,-94</points>
<intersection>19 0</intersection>
<intersection>71 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>71,-94,71,-19.5</points>
<intersection>-94 2</intersection>
<intersection>-19.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>63.5,-19.5,72,-19.5</points>
<connection>
<GID>93</GID>
<name>OUT_0</name></connection>
<connection>
<GID>110</GID>
<name>N_in0</name></connection>
<intersection>71 3</intersection></hsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-93,20,-46.5</points>
<intersection>-93 1</intersection>
<intersection>-46.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20,-93,70,-93</points>
<intersection>20 0</intersection>
<intersection>70 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>20,-46.5,27,-46.5</points>
<connection>
<GID>97</GID>
<name>IN_1</name></connection>
<intersection>20 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>70,-93,70,-28</points>
<intersection>-93 1</intersection>
<intersection>-28 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>63.5,-28,72,-28</points>
<connection>
<GID>94</GID>
<name>OUT_0</name></connection>
<connection>
<GID>111</GID>
<name>N_in0</name></connection>
<intersection>70 3</intersection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-92,69,-36.5</points>
<intersection>-92 1</intersection>
<intersection>-36.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,-92,69,-92</points>
<intersection>21 3</intersection>
<intersection>69 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,-36.5,72,-36.5</points>
<connection>
<GID>95</GID>
<name>OUT_0</name></connection>
<connection>
<GID>112</GID>
<name>N_in0</name></connection>
<intersection>69 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>21,-92,21,-47.5</points>
<intersection>-92 1</intersection>
<intersection>-47.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>21,-47.5,27,-47.5</points>
<connection>
<GID>97</GID>
<name>IN_2</name></connection>
<intersection>21 3</intersection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-91,22,-48.5</points>
<intersection>-91 2</intersection>
<intersection>-48.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22,-48.5,27,-48.5</points>
<connection>
<GID>97</GID>
<name>IN_3</name></connection>
<intersection>22 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-91,68,-91</points>
<intersection>22 0</intersection>
<intersection>68 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>68,-91,68,-45</points>
<intersection>-91 2</intersection>
<intersection>-45 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>63.5,-45,72,-45</points>
<connection>
<GID>96</GID>
<name>OUT_0</name></connection>
<connection>
<GID>113</GID>
<name>N_in0</name></connection>
<intersection>68 3</intersection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-90,23,-62.5</points>
<intersection>-90 2</intersection>
<intersection>-62.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-62.5,27,-62.5</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23,-90,67,-90</points>
<intersection>23 0</intersection>
<intersection>67 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>67,-90,67,-55</points>
<intersection>-90 2</intersection>
<intersection>-55 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>63.5,-55,72,-55</points>
<connection>
<GID>106</GID>
<name>OUT_0</name></connection>
<connection>
<GID>114</GID>
<name>N_in0</name></connection>
<intersection>67 3</intersection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24,-89,66,-89</points>
<intersection>24 3</intersection>
<intersection>66 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>24,-89,24,-63.5</points>
<intersection>-89 1</intersection>
<intersection>-63.5 5</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>66,-89,66,-63.5</points>
<intersection>-89 1</intersection>
<intersection>-63.5 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>24,-63.5,27,-63.5</points>
<connection>
<GID>101</GID>
<name>IN_1</name></connection>
<intersection>24 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>63.5,-63.5,72,-63.5</points>
<connection>
<GID>107</GID>
<name>OUT_0</name></connection>
<connection>
<GID>115</GID>
<name>N_in0</name></connection>
<intersection>66 4</intersection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,-88,65,-72</points>
<intersection>-88 1</intersection>
<intersection>-72 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-88,65,-88</points>
<intersection>25 3</intersection>
<intersection>65 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,-72,72,-72</points>
<connection>
<GID>108</GID>
<name>OUT_0</name></connection>
<connection>
<GID>116</GID>
<name>N_in0</name></connection>
<intersection>65 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>25,-88,25,-64.5</points>
<intersection>-88 1</intersection>
<intersection>-64.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>25,-64.5,27,-64.5</points>
<connection>
<GID>101</GID>
<name>IN_2</name></connection>
<intersection>25 3</intersection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,-87,64,-80.5</points>
<intersection>-87 1</intersection>
<intersection>-80.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-87,64,-87</points>
<intersection>26 3</intersection>
<intersection>64 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,-80.5,72.5,-80.5</points>
<connection>
<GID>109</GID>
<name>OUT_0</name></connection>
<connection>
<GID>117</GID>
<name>N_in0</name></connection>
<intersection>64 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>26,-87,26,-65.5</points>
<intersection>-87 1</intersection>
<intersection>-65.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>26,-65.5,27,-65.5</points>
<connection>
<GID>101</GID>
<name>IN_3</name></connection>
<intersection>26 3</intersection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,-80.5,95,-80.5</points>
<connection>
<GID>117</GID>
<name>N_in1</name></connection>
<connection>
<GID>118</GID>
<name>ADDRESS_7</name></connection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-81.5,76,-72</points>
<intersection>-81.5 2</intersection>
<intersection>-72 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74,-72,76,-72</points>
<connection>
<GID>116</GID>
<name>N_in1</name></connection>
<intersection>76 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>76,-81.5,95,-81.5</points>
<connection>
<GID>118</GID>
<name>ADDRESS_6</name></connection>
<intersection>76 0</intersection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77,-82.5,77,-63.5</points>
<intersection>-82.5 2</intersection>
<intersection>-63.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74,-63.5,77,-63.5</points>
<connection>
<GID>115</GID>
<name>N_in1</name></connection>
<intersection>77 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77,-82.5,95,-82.5</points>
<connection>
<GID>118</GID>
<name>ADDRESS_5</name></connection>
<intersection>77 0</intersection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78,-83.5,78,-55</points>
<intersection>-83.5 2</intersection>
<intersection>-55 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74,-55,78,-55</points>
<connection>
<GID>114</GID>
<name>N_in1</name></connection>
<intersection>78 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>78,-83.5,95,-83.5</points>
<connection>
<GID>118</GID>
<name>ADDRESS_4</name></connection>
<intersection>78 0</intersection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79,-84.5,79,-45</points>
<intersection>-84.5 2</intersection>
<intersection>-45 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74,-45,79,-45</points>
<connection>
<GID>113</GID>
<name>N_in1</name></connection>
<intersection>79 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>79,-84.5,95,-84.5</points>
<connection>
<GID>118</GID>
<name>ADDRESS_3</name></connection>
<intersection>79 0</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-85.5,80,-36.5</points>
<intersection>-85.5 2</intersection>
<intersection>-36.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74,-36.5,80,-36.5</points>
<connection>
<GID>112</GID>
<name>N_in1</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>80,-85.5,95,-85.5</points>
<connection>
<GID>118</GID>
<name>ADDRESS_2</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,-86.5,81,-28</points>
<intersection>-86.5 2</intersection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74,-28,81,-28</points>
<connection>
<GID>111</GID>
<name>N_in1</name></connection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>81,-86.5,95,-86.5</points>
<connection>
<GID>118</GID>
<name>ADDRESS_1</name></connection>
<intersection>81 0</intersection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82,-87.5,82,-19.5</points>
<intersection>-87.5 2</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74,-19.5,82,-19.5</points>
<connection>
<GID>110</GID>
<name>N_in1</name></connection>
<intersection>82 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>82,-87.5,95,-87.5</points>
<connection>
<GID>118</GID>
<name>ADDRESS_0</name></connection>
<intersection>82 0</intersection></hsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>105,-84.5,106,-84.5</points>
<connection>
<GID>118</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>119</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,38.5,22,39.5</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>38.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,38.5,55,38.5</points>
<connection>
<GID>124</GID>
<name>N_in1</name></connection>
<intersection>22 0</intersection>
<intersection>55 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>55,38.5,55,55.5</points>
<connection>
<GID>147</GID>
<name>IN_0</name></connection>
<intersection>38.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21,37.5,62,37.5</points>
<connection>
<GID>125</GID>
<name>N_in1</name></connection>
<intersection>26 2</intersection>
<intersection>62 4</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>26,37.5,26,39.5</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<intersection>37.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>62,37.5,62,55.5</points>
<connection>
<GID>149</GID>
<name>IN_1</name></connection>
<intersection>37.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,36.5,30,39.5</points>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<intersection>36.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,36.5,71,36.5</points>
<connection>
<GID>126</GID>
<name>N_in1</name></connection>
<intersection>30 0</intersection>
<intersection>71 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>71,36.5,71,55.5</points>
<connection>
<GID>151</GID>
<name>IN_2</name></connection>
<intersection>36.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,35.5,34,39.5</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<intersection>35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,35.5,86,35.5</points>
<connection>
<GID>127</GID>
<name>N_in1</name></connection>
<intersection>34 0</intersection>
<intersection>86 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>86,35.5,86,55.5</points>
<connection>
<GID>154</GID>
<name>IN_1</name></connection>
<intersection>35.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,34.5,38,39.5</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<intersection>34.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,34.5,103,34.5</points>
<connection>
<GID>128</GID>
<name>N_in1</name></connection>
<intersection>38 0</intersection>
<intersection>103 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>103,34.5,103,55.5</points>
<connection>
<GID>157</GID>
<name>IN_1</name></connection>
<intersection>34.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,32.5,46,39.5</points>
<connection>
<GID>134</GID>
<name>IN_0</name></connection>
<intersection>32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,32.5,132.5,32.5</points>
<connection>
<GID>130</GID>
<name>N_in1</name></connection>
<intersection>46 0</intersection>
<intersection>132.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>132.5,32.5,132.5,55.5</points>
<connection>
<GID>165</GID>
<name>IN_6</name></connection>
<intersection>32.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,31.5,50,39.5</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<intersection>31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,31.5,142.5,31.5</points>
<connection>
<GID>131</GID>
<name>N_in1</name></connection>
<intersection>50 0</intersection>
<intersection>142.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>142.5,31.5,142.5,55.5</points>
<connection>
<GID>161</GID>
<name>IN_7</name></connection>
<intersection>31.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,26.5,24,39.5</points>
<connection>
<GID>120</GID>
<name>IN_1</name></connection>
<intersection>26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,26.5,57,26.5</points>
<connection>
<GID>136</GID>
<name>N_in1</name></connection>
<intersection>24 0</intersection>
<intersection>57 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>57,26.5,57,39.5</points>
<connection>
<GID>148</GID>
<name>IN_0</name></connection>
<intersection>26.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,25.5,28,39.5</points>
<connection>
<GID>121</GID>
<name>IN_1</name></connection>
<intersection>25.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,25.5,64,25.5</points>
<connection>
<GID>137</GID>
<name>N_in1</name></connection>
<intersection>28 0</intersection>
<intersection>64 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>64,25.5,64,39.5</points>
<connection>
<GID>150</GID>
<name>IN_0</name></connection>
<intersection>25.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,24.5,32,39.5</points>
<connection>
<GID>122</GID>
<name>IN_1</name></connection>
<intersection>24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,24.5,73,24.5</points>
<connection>
<GID>138</GID>
<name>N_in1</name></connection>
<intersection>32 0</intersection>
<intersection>73 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>73,24.5,73,39.5</points>
<connection>
<GID>152</GID>
<name>IN_0</name></connection>
<intersection>24.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,23.5,36,39.5</points>
<connection>
<GID>123</GID>
<name>IN_1</name></connection>
<intersection>23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,23.5,88,23.5</points>
<connection>
<GID>139</GID>
<name>N_in1</name></connection>
<intersection>36 0</intersection>
<intersection>88 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>88,23.5,88,39.5</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<intersection>23.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,22.5,40,39.5</points>
<connection>
<GID>132</GID>
<name>IN_1</name></connection>
<intersection>22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,22.5,105,22.5</points>
<connection>
<GID>140</GID>
<name>N_in1</name></connection>
<intersection>40 0</intersection>
<intersection>105 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>105,22.5,105,39.5</points>
<connection>
<GID>158</GID>
<name>IN_0</name></connection>
<intersection>22.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,21.5,44,39.5</points>
<connection>
<GID>133</GID>
<name>IN_1</name></connection>
<intersection>21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,21.5,124,21.5</points>
<connection>
<GID>141</GID>
<name>N_in1</name></connection>
<intersection>44 0</intersection>
<intersection>124 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>124,21.5,124,39.5</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<intersection>21.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48,20.5,48,39.5</points>
<connection>
<GID>134</GID>
<name>IN_1</name></connection>
<intersection>20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,20.5,133.5,20.5</points>
<connection>
<GID>142</GID>
<name>N_in1</name></connection>
<intersection>48 0</intersection>
<intersection>133.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>133.5,20.5,133.5,39.5</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>20.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,19.5,52,39.5</points>
<connection>
<GID>135</GID>
<name>IN_1</name></connection>
<intersection>19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,19.5,148,19.5</points>
<connection>
<GID>143</GID>
<name>N_in1</name></connection>
<intersection>52 0</intersection>
<intersection>148 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>148,19.5,148,39.5</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<intersection>19.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>27,45.5,27,47.5</points>
<connection>
<GID>121</GID>
<name>OUT</name></connection>
<intersection>47.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>9,47.5,136.5,47.5</points>
<intersection>9 3</intersection>
<intersection>27 1</intersection>
<intersection>69 5</intersection>
<intersection>78 7</intersection>
<intersection>93 9</intersection>
<intersection>110 12</intersection>
<intersection>127.5 15</intersection>
<intersection>136.5 14</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>9,47.5,9,54.5</points>
<connection>
<GID>144</GID>
<name>IN_1</name></connection>
<intersection>47.5 2</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>69,47.5,69,55.5</points>
<connection>
<GID>151</GID>
<name>IN_1</name></connection>
<intersection>47.5 2</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>78,47.5,78,55.5</points>
<connection>
<GID>153</GID>
<name>IN_1</name></connection>
<intersection>47.5 2</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>93,47.5,93,55.5</points>
<connection>
<GID>156</GID>
<name>IN_1</name></connection>
<intersection>47.5 2</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>110,47.5,110,55.5</points>
<connection>
<GID>159</GID>
<name>IN_1</name></connection>
<intersection>47.5 2</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>136.5,47.5,136.5,55.5</points>
<connection>
<GID>161</GID>
<name>IN_1</name></connection>
<intersection>47.5 2</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>127.5,47.5,127.5,55.5</points>
<connection>
<GID>165</GID>
<name>IN_1</name></connection>
<intersection>47.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,48.5,11,54.5</points>
<connection>
<GID>144</GID>
<name>IN_2</name></connection>
<intersection>48.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>31,45.5,31,48.5</points>
<connection>
<GID>122</GID>
<name>OUT</name></connection>
<intersection>48.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>11,48.5,137.5,48.5</points>
<intersection>11 0</intersection>
<intersection>31 1</intersection>
<intersection>80 4</intersection>
<intersection>95 6</intersection>
<intersection>112 9</intersection>
<intersection>128.5 12</intersection>
<intersection>137.5 11</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>80,48.5,80,55.5</points>
<connection>
<GID>153</GID>
<name>IN_2</name></connection>
<intersection>48.5 2</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>95,48.5,95,55.5</points>
<connection>
<GID>156</GID>
<name>IN_2</name></connection>
<intersection>48.5 2</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>112,48.5,112,55.5</points>
<connection>
<GID>159</GID>
<name>IN_2</name></connection>
<intersection>48.5 2</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>137.5,48.5,137.5,55.5</points>
<connection>
<GID>161</GID>
<name>IN_2</name></connection>
<intersection>48.5 2</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>128.5,48.5,128.5,55.5</points>
<connection>
<GID>165</GID>
<name>IN_2</name></connection>
<intersection>48.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,46.5,7,54.5</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<intersection>46.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>7,46.5,135.5,46.5</points>
<intersection>7 0</intersection>
<intersection>23 4</intersection>
<intersection>60 5</intersection>
<intersection>67 7</intersection>
<intersection>76 9</intersection>
<intersection>91 11</intersection>
<intersection>108 14</intersection>
<intersection>126.5 17</intersection>
<intersection>135.5 16</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>23,45.5,23,46.5</points>
<connection>
<GID>120</GID>
<name>OUT</name></connection>
<intersection>46.5 3</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>60,46.5,60,55.5</points>
<connection>
<GID>149</GID>
<name>IN_0</name></connection>
<intersection>46.5 3</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>67,46.5,67,55.5</points>
<connection>
<GID>151</GID>
<name>IN_0</name></connection>
<intersection>46.5 3</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>76,46.5,76,55.5</points>
<connection>
<GID>153</GID>
<name>IN_0</name></connection>
<intersection>46.5 3</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>91,46.5,91,55.5</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<intersection>46.5 3</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>108,46.5,108,55.5</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<intersection>46.5 3</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>135.5,46.5,135.5,55.5</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<intersection>46.5 3</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>126.5,46.5,126.5,55.5</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<intersection>46.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,45.5,35,49.5</points>
<connection>
<GID>123</GID>
<name>OUT</name></connection>
<intersection>49.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>13,49.5,13,54.5</points>
<connection>
<GID>144</GID>
<name>IN_3</name></connection>
<intersection>49.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>13,49.5,138.5,49.5</points>
<intersection>13 1</intersection>
<intersection>35 0</intersection>
<intersection>97 4</intersection>
<intersection>114 6</intersection>
<intersection>129.5 9</intersection>
<intersection>138.5 8</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>97,49.5,97,55.5</points>
<connection>
<GID>156</GID>
<name>IN_3</name></connection>
<intersection>49.5 2</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>114,49.5,114,55.5</points>
<connection>
<GID>159</GID>
<name>IN_3</name></connection>
<intersection>49.5 2</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>138.5,49.5,138.5,55.5</points>
<connection>
<GID>161</GID>
<name>IN_3</name></connection>
<intersection>49.5 2</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>129.5,49.5,129.5,55.5</points>
<connection>
<GID>165</GID>
<name>IN_3</name></connection>
<intersection>49.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,45.5,43,51.5</points>
<connection>
<GID>133</GID>
<name>OUT</name></connection>
<intersection>51.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>17,51.5,17,54.5</points>
<connection>
<GID>145</GID>
<name>IN_1</name></connection>
<intersection>51.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>17,51.5,140.5,51.5</points>
<intersection>17 1</intersection>
<intersection>43 0</intersection>
<intersection>131.5 7</intersection>
<intersection>140.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>140.5,51.5,140.5,55.5</points>
<connection>
<GID>161</GID>
<name>IN_5</name></connection>
<intersection>51.5 2</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>131.5,51.5,131.5,55.5</points>
<connection>
<GID>165</GID>
<name>IN_5</name></connection>
<intersection>51.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,45.5,47,52.5</points>
<connection>
<GID>134</GID>
<name>OUT</name></connection>
<intersection>52.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>19,52.5,19,54.5</points>
<connection>
<GID>145</GID>
<name>IN_2</name></connection>
<intersection>52.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>19,52.5,141.5,52.5</points>
<intersection>19 1</intersection>
<intersection>47 0</intersection>
<intersection>141.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>141.5,52.5,141.5,55.5</points>
<connection>
<GID>161</GID>
<name>IN_6</name></connection>
<intersection>52.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,45.5,39,50.5</points>
<connection>
<GID>132</GID>
<name>OUT</name></connection>
<intersection>50.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>15,50.5,15,54.5</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<intersection>50.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>15,50.5,139.5,50.5</points>
<intersection>15 1</intersection>
<intersection>39 0</intersection>
<intersection>120 6</intersection>
<intersection>130.5 9</intersection>
<intersection>139.5 8</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>120,50.5,120,55.5</points>
<connection>
<GID>160</GID>
<name>IN_1</name></connection>
<intersection>50.5 2</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>139.5,50.5,139.5,55.5</points>
<connection>
<GID>161</GID>
<name>IN_4</name></connection>
<intersection>50.5 2</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>130.5,50.5,130.5,55.5</points>
<connection>
<GID>165</GID>
<name>IN_4</name></connection>
<intersection>50.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>10,61.5,13,61.5</points>
<intersection>10 4</intersection>
<intersection>13 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>13,61.5,13,62.5</points>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<intersection>61.5 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>10,60.5,10,61.5</points>
<connection>
<GID>144</GID>
<name>OUT</name></connection>
<intersection>61.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,60.5,18,61.5</points>
<connection>
<GID>145</GID>
<name>OUT</name></connection>
<intersection>61.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>15,61.5,15,62.5</points>
<connection>
<GID>146</GID>
<name>IN_1</name></connection>
<intersection>61.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>15,61.5,18,61.5</points>
<intersection>15 1</intersection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,43.5,57,55.5</points>
<connection>
<GID>148</GID>
<name>OUT_0</name></connection>
<connection>
<GID>147</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,43.5,64,55.5</points>
<connection>
<GID>150</GID>
<name>OUT_0</name></connection>
<connection>
<GID>149</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,43.5,73,55.5</points>
<connection>
<GID>152</GID>
<name>OUT_0</name></connection>
<connection>
<GID>151</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82,54.5,82,62.5</points>
<intersection>54.5 4</intersection>
<intersection>62.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>78,62.5,82,62.5</points>
<intersection>78 7</intersection>
<intersection>82 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>82,54.5,84,54.5</points>
<intersection>82 0</intersection>
<intersection>84 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>84,54.5,84,55.5</points>
<connection>
<GID>154</GID>
<name>IN_0</name></connection>
<intersection>54.5 4</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>78,61.5,78,62.5</points>
<connection>
<GID>153</GID>
<name>OUT</name></connection>
<intersection>62.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,43.5,88,55.5</points>
<connection>
<GID>155</GID>
<name>OUT_0</name></connection>
<connection>
<GID>154</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,54.5,99,62.5</points>
<intersection>54.5 3</intersection>
<intersection>62.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>94,61.5,94,62.5</points>
<connection>
<GID>156</GID>
<name>OUT</name></connection>
<intersection>62.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>94,62.5,99,62.5</points>
<intersection>94 1</intersection>
<intersection>99 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>99,54.5,101,54.5</points>
<intersection>99 0</intersection>
<intersection>101 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>101,54.5,101,55.5</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>54.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105,43.5,105,55.5</points>
<connection>
<GID>158</GID>
<name>OUT_0</name></connection>
<connection>
<GID>157</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,33.5,42,39.5</points>
<connection>
<GID>133</GID>
<name>IN_0</name></connection>
<intersection>33.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,33.5,122,33.5</points>
<connection>
<GID>129</GID>
<name>N_in1</name></connection>
<intersection>42 0</intersection>
<intersection>122 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>122,33.5,122,55.5</points>
<connection>
<GID>160</GID>
<name>IN_2</name></connection>
<intersection>33.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,61.5,111,62.5</points>
<connection>
<GID>159</GID>
<name>OUT</name></connection>
<intersection>62.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>116,54.5,116,62.5</points>
<intersection>54.5 3</intersection>
<intersection>62.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>111,62.5,116,62.5</points>
<intersection>111 0</intersection>
<intersection>116 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>116,54.5,118,54.5</points>
<intersection>116 1</intersection>
<intersection>118 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>118,54.5,118,55.5</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<intersection>54.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21,53.5,21,54.5</points>
<connection>
<GID>145</GID>
<name>IN_3</name></connection>
<intersection>53.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>51,45.5,51,53.5</points>
<connection>
<GID>135</GID>
<name>OUT</name></connection>
<intersection>53.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>21,53.5,51,53.5</points>
<intersection>21 0</intersection>
<intersection>51 1</intersection></hsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139,61.5,139,62.5</points>
<connection>
<GID>161</GID>
<name>OUT</name></connection>
<intersection>62.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>144,55.5,144,62.5</points>
<intersection>55.5 3</intersection>
<intersection>62.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>139,62.5,144,62.5</points>
<intersection>139 0</intersection>
<intersection>144 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>144,55.5,146,55.5</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<intersection>144 1</intersection></hsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148,43.5,148,55.5</points>
<connection>
<GID>163</GID>
<name>OUT_0</name></connection>
<connection>
<GID>162</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124,43.5,124,55.5</points>
<connection>
<GID>164</GID>
<name>OUT_0</name></connection>
<connection>
<GID>160</GID>
<name>IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133.5,43.5,133.5,55.5</points>
<connection>
<GID>166</GID>
<name>OUT_0</name></connection>
<connection>
<GID>165</GID>
<name>IN_7</name></connection></vsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,62.5,46.5,70.5</points>
<connection>
<GID>167</GID>
<name>IN_0</name></connection>
<intersection>62.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>56,61.5,56,62.5</points>
<connection>
<GID>147</GID>
<name>OUT</name></connection>
<intersection>62.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>46.5,62.5,56,62.5</points>
<intersection>46.5 0</intersection>
<intersection>56 1</intersection></hsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,63.5,47.5,70.5</points>
<connection>
<GID>167</GID>
<name>IN_1</name></connection>
<intersection>63.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>62,61.5,62,63.5</points>
<connection>
<GID>149</GID>
<name>OUT</name></connection>
<intersection>63.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>47.5,63.5,62,63.5</points>
<intersection>47.5 0</intersection>
<intersection>62 1</intersection></hsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48.5,64.5,48.5,70.5</points>
<connection>
<GID>167</GID>
<name>IN_2</name></connection>
<intersection>64.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>70,61.5,70,64.5</points>
<connection>
<GID>151</GID>
<name>OUT</name></connection>
<intersection>64.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>48.5,64.5,70,64.5</points>
<intersection>48.5 0</intersection>
<intersection>70 1</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>0,492.194,1138,-368.806</PageViewport></page 2>
<page 3>
<PageViewport>0,492.194,1138,-368.806</PageViewport></page 3>
<page 4>
<PageViewport>0,492.194,1138,-368.806</PageViewport></page 4>
<page 5>
<PageViewport>0,492.194,1138,-368.806</PageViewport></page 5>
<page 6>
<PageViewport>0,492.194,1138,-368.806</PageViewport></page 6>
<page 7>
<PageViewport>0,492.194,1138,-368.806</PageViewport></page 7>
<page 8>
<PageViewport>0,492.194,1138,-368.806</PageViewport></page 8>
<page 9>
<PageViewport>0,492.194,1138,-368.806</PageViewport></page 9></circuit>